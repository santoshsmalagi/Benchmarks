//# 28 inputs
//# 106 outputs
//# 1636 D-type flipflops
//# 13470 inverters
//# 8709 gates (4154 ANDs + 2050 NANDs + 226 ORs + 2279 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;
reg Q;
always @ (posedge CK)
  Q <= D;
endmodule

module s38417(CK,g1249,g16297,g16355,g16399,g16437,g16496,g1943,g24734,
  g25420,
  g25435,g25442,g25489,g26104,g26135,g26149,g2637,g27380,g3212,g3213,g3214,
  g3215,g3216,g3217,g3218,g3219,g3220,g3221,g3222,g3223,g3224,g3225,g3226,
  g3227,g3228,g3229,g3230,g3231,g3232,g3233,g3234,g3993,g4088,g4090,g4200,
  g4321,g4323,g4450,g4590,g51,g5388,g5437,g5472,g5511,g5549,g5555,g5595,g5612,
  g5629,g563,g5637,g5648,g5657,g5686,g5695,g5738,g5747,g5796,g6225,g6231,g6313,
  g6368,g6442,g6447,g6485,g6518,g6573,g6642,g6677,g6712,g6750,g6782,g6837,
  g6895,g6911,g6944,g6979,g7014,g7052,g7084,g7161,g7194,g7229,g7264,g7302,
  g7334,g7357,g7390,g7425,g7487,g7519,g7909,g7956,g7961,g8007,g8012,g8021,
  g8023,g8030,g8082,g8087,g8096,g8106,g8167,g8175,g8249,g8251,g8258,g8259,
  g8260,g8261,g8262,g8263,g8264,g8265,g8266,g8267,g8268,g8269,g8270,g8271,
  g8272,g8273,g8274,g8275);
input CK,g51,g563,g1249,g1943,g2637,g3212,g3213,g3214,g3215,g3216,
  g3217,g3218,
  g3219,g3220,g3221,g3222,g3223,g3224,g3225,g3226,g3227,g3228,g3229,g3230,
  g3231,g3232,g3233,g3234;
output g3993,g4088,g4090,g4200,g4321,g4323,g4450,g4590,g5388,g5437,g5472,g5511,
  g5549,g5555,g5595,g5612,g5629,g5637,g5648,g5657,g5686,g5695,g5738,g5747,
  g5796,g6225,g6231,g6313,g6368,g6442,g6447,g6485,g6518,g6573,g6642,g6677,
  g6712,g6750,g6782,g6837,g6895,g6911,g6944,g6979,g7014,g7052,g7084,g7161,
  g7194,g7229,g7264,g7302,g7334,g7357,g7390,g7425,g7487,g7519,g7909,g7956,
  g7961,g8007,g8012,g8021,g8023,g8030,g8082,g8087,g8096,g8106,g8167,g8175,
  g8249,g8251,g8258,g8259,g8260,g8261,g8262,g8263,g8264,g8265,g8266,g8267,
  g8268,g8269,g8270,g8271,g8272,g8273,g8274,g8275,g16297,g16355,g16399,g16437,
  g16496,g24734,g25420,g25435,g25442,g25489,g26104,g26135,g26149,g27380;

  wire g2814,g16475,g2817,g20571,g2933,g20588,g2950,g21951,g2883,g23315,g2888,
    g24423,g2896,g25175,g2892,g26019,g2903,g26747,g2900,g27237,g2908,g27715,
    g2912,g24424,g2917,g25174,g2924,g26020,g2920,g26746,g2984,g19061,g2985,
    g19060,g2930,g19062,g2929,g2879,g16494,g2934,g16476,g2935,g16477,g2938,
    g16478,g2941,g16479,g2944,g16480,g2947,g16481,g2953,g16482,g2956,g16483,
    g2959,g16484,g2962,g16485,g2963,g16486,g2966,g16487,g2969,g16488,g2972,
    g16489,g2975,g16490,g2978,g16491,g2981,g16492,g2874,g16493,g1506,g20572,
    g1501,g20573,g1496,g20574,g1491,g20575,g1486,g20576,g1481,g20577,g1476,
    g20578,g1471,g20579,g2877,g23313,g2861,g21960,g813,g2864,g21961,g809,g2867,
    g21962,g805,g2870,g21963,g801,g2818,g21947,g797,g2821,g21948,g793,g2824,
    g21949,g789,g2827,g21950,g785,g2830,g23312,g2873,g2833,g21952,g125,g2836,
    g21953,g121,g2839,g21954,g117,g2842,g21955,g113,g2845,g21956,g109,g2848,
    g21957,g105,g2851,g21958,g101,g2854,g21959,g97,g2858,g23316,g2857,g2200,
    g20587,g2195,g20585,g2190,g20586,g2185,g20584,g2180,g20583,g2175,g20582,
    g2170,g20581,g2165,g20580,g2878,g23314,g3129,g13475,g3117,g3109,g3210,
    g20630,g3211,g20631,g3084,g20632,g3085,g20609,g3086,g20610,g3087,g20611,
    g3091,g20612,g3092,g20613,g3093,g20614,g3094,g20615,g3095,g20616,g3096,
    g20617,g3097,g26751,g3098,g26752,g3099,g26753,g3100,g29163,g3101,g29164,
    g3102,g29165,g3103,g30120,g3104,g30121,g3105,g30122,g3106,g30941,g3107,
    g30942,g3108,g30943,g3155,g20618,g3158,g20619,g3161,g20620,g3164,g20621,
    g3167,g20622,g3170,g20623,g3173,g20624,g3176,g20625,g3179,g20626,g3182,
    g20627,g3185,g20628,g3088,g20629,g3191,g27717,g3194,g28316,g3197,g28317,
    g3198,g28318,g3201,g28704,g3204,g28705,g3207,g28706,g3188,g29463,g3133,
    g29656,g3132,g28698,g3128,g29166,g3127,g28697,g3126,g28315,g3125,g28696,
    g3124,g28314,g3123,g28313,g3120,g28695,g3114,g28694,g3113,g28693,g3112,
    g28312,g3110,g28311,g3111,g28310,g3139,g29461,g3136,g28701,g3134,g28700,
    g3135,g28699,g3151,g29462,g3142,g28703,g3147,g28702,g185,g29657,g138,
    g13405,g135,g165,g130,g24259,g131,g24260,g129,g24261,g133,g24262,g134,
    g24263,g132,g24264,g142,g24265,g143,g24266,g141,g24267,g145,g24268,g146,
    g24269,g144,g24270,g148,g24271,g149,g24272,g147,g24273,g151,g24274,g152,
    g24275,g150,g24276,g154,g24277,g155,g24278,g153,g24279,g157,g24280,g158,
    g24281,g156,g24282,g160,g24283,g161,g24284,g159,g24285,g163,g24286,g164,
    g24287,g162,g24288,g169,g26679,g170,g26680,g168,g26681,g172,g26682,g173,
    g26683,g171,g26684,g175,g26685,g176,g26686,g174,g26687,g178,g26688,g179,
    g26689,g177,g26690,g186,g30506,g189,g30507,g192,g30508,g231,g30842,g234,
    g30843,g237,g30844,g195,g30836,g198,g30837,g201,g30838,g240,g30845,g243,
    g30846,g246,g30847,g204,g30509,g207,g30510,g210,g30511,g249,g30515,g252,
    g30516,g255,g30517,g213,g30512,g216,g30513,g219,g30514,g258,g30518,g261,
    g30519,g264,g30520,g222,g30839,g225,g30840,g228,g30841,g267,g30848,g270,
    g30849,g273,g30850,g92,g25983,g88,g26678,g83,g27189,g79,g27683,g74,g28206,
    g70,g28673,g65,g29131,g61,g29413,g56,g29627,g52,g29794,g180,g20555,g182,
    g181,g276,g13406,g405,g401,g309,g11496,g354,g28207,g343,g28208,g346,g28209,
    g369,g28210,g358,g28211,g361,g28212,g384,g28213,g373,g28214,g376,g28215,
    g398,g28216,g388,g28217,g391,g28218,g408,g29414,g411,g29415,g414,g29416,
    g417,g29631,g420,g29632,g423,g29633,g427,g29417,g428,g29418,g426,g29419,
    g429,g27684,g432,g27685,g435,g27686,g438,g27687,g441,g27688,g444,g27689,
    g448,g28674,g449,g28675,g447,g28676,g312,g29795,g313,g29796,g314,g29797,
    g315,g30851,g316,g30852,g317,g30853,g318,g30710,g319,g30711,g320,g30712,
    g322,g29628,g323,g29629,g321,g29630,g403,g27191,g404,g27192,g402,g27193,
    g450,g11509,g451,g452,g11510,g453,g454,g11511,g279,g280,g11491,g281,g282,
    g11492,g283,g284,g11493,g285,g286,g11494,g287,g288,g11495,g289,g290,g13407,
    g291,g299,g19012,g305,g23148,g308,g23149,g297,g23150,g296,g23151,g295,
    g23152,g294,g23153,g304,g19016,g303,g19015,g302,g19014,g301,g19013,g300,
    g25130,g298,g27190,g342,g11497,g349,g350,g11498,g351,g352,g11499,g353,g357,
    g11500,g364,g365,g11501,g366,g367,g11502,g368,g372,g11503,g379,g380,g11504,
    g381,g382,g11505,g383,g387,g11506,g394,g395,g11507,g396,g397,g11508,g324,
    g325,g13408,g331,g337,g545,g13419,g551,g550,g554,g23160,g557,g20556,g510,
    g20557,g513,g16467,g523,g524,g564,g11512,g569,g570,g11515,g571,g572,g11516,
    g573,g574,g11517,g565,g566,g11513,g567,g568,g11514,g489,g474,g13409,g481,
    g485,g486,g24292,g487,g24293,g488,g24294,g455,g25139,g458,g25131,g461,
    g25132,g477,g25136,g478,g25137,g479,g25138,g480,g24289,g484,g24290,g464,
    g24291,g465,g25133,g468,g25134,g471,g25135,g528,g16468,g535,g542,g543,
    g19021,g544,g548,g23159,g549,g19022,g499,g558,g19023,g559,g576,g28219,g577,
    g28220,g575,g28221,g579,g28222,g580,g28223,g578,g28224,g582,g28225,g583,
    g28226,g581,g28227,g585,g28228,g586,g28229,g584,g28230,g587,g25985,g590,
    g25986,g593,g25987,g596,g25988,g599,g25989,g602,g25990,g614,g29135,g617,
    g29136,g620,g29137,g605,g29132,g608,g29133,g611,g29134,g490,g27194,g493,
    g27195,g496,g27196,g506,g8284,g507,g24295,g508,g19017,g509,g19018,g514,
    g19019,g515,g19020,g516,g23158,g517,g23157,g518,g23156,g519,g23155,g520,
    g23154,g525,g529,g13410,g530,g13411,g531,g13412,g532,g13413,g533,g13414,
    g534,g13415,g536,g13416,g537,g13417,g538,g25984,g541,g13418,g623,g13420,
    g626,g629,g630,g20558,g659,g21943,g640,g23161,g633,g24296,g653,g25140,g646,
    g25991,g660,g26691,g672,g27197,g666,g27690,g679,g28231,g686,g28677,g692,
    g29138,g699,g23162,g700,g23163,g698,g23164,g702,g23165,g703,g23166,g701,
    g23167,g705,g23168,g706,g23169,g704,g23170,g708,g23171,g709,g23172,g707,
    g23173,g711,g23174,g712,g23175,g710,g23176,g714,g23177,g715,g23178,g713,
    g23179,g717,g23180,g718,g23181,g716,g23182,g720,g23183,g721,g23184,g719,
    g23185,g723,g23186,g724,g23187,g722,g23188,g726,g23189,g727,g23190,g725,
    g23191,g729,g23192,g730,g23193,g728,g23194,g732,g23195,g733,g23196,g731,
    g23197,g735,g26692,g736,g26693,g734,g26694,g738,g24297,g739,g24298,g737,
    g24299,g826,g13421,g823,g853,g818,g24300,g819,g24301,g817,g24302,g821,
    g24303,g822,g24304,g820,g24305,g830,g24306,g831,g24307,g829,g24308,g833,
    g24309,g834,g24310,g832,g24311,g836,g24312,g837,g24313,g835,g24314,g839,
    g24315,g840,g24316,g838,g24317,g842,g24318,g843,g24319,g841,g24320,g845,
    g24321,g846,g24322,g844,g24323,g848,g24324,g849,g24325,g847,g24326,g851,
    g24327,g852,g24328,g850,g24329,g857,g26696,g858,g26697,g856,g26698,g860,
    g26699,g861,g26700,g859,g26701,g863,g26702,g864,g26703,g862,g26704,g866,
    g26705,g867,g26706,g865,g26707,g873,g30521,g876,g30522,g879,g30523,g918,
    g30860,g921,g30861,g924,g30862,g882,g30854,g885,g30855,g888,g30856,g927,
    g30863,g930,g30864,g933,g30865,g891,g30524,g894,g30525,g897,g30526,g936,
    g30530,g939,g30531,g942,g30532,g900,g30527,g903,g30528,g906,g30529,g945,
    g30533,g948,g30534,g951,g30535,g909,g30857,g912,g30858,g915,g30859,g954,
    g30866,g957,g30867,g960,g30868,g780,g25992,g776,g26695,g771,g27198,g767,
    g27691,g762,g28232,g758,g28678,g753,g29139,g749,g29420,g744,g29634,g740,
    g29798,g868,g20559,g870,g869,g963,g13422,g1092,g1088,g996,g11523,g1041,
    g28233,g1030,g28234,g1033,g28235,g1056,g28236,g1045,g28237,g1048,g28238,
    g1071,g28239,g1060,g28240,g1063,g28241,g1085,g28242,g1075,g28243,g1078,
    g28244,g1095,g29421,g1098,g29422,g1101,g29423,g1104,g29638,g1107,g29639,
    g1110,g29640,g1114,g29424,g1115,g29425,g1113,g29426,g1116,g27692,g1119,
    g27693,g1122,g27694,g1125,g27695,g1128,g27696,g1131,g27697,g1135,g28679,
    g1136,g28680,g1134,g28681,g999,g29799,g1000,g29800,g1001,g29801,g1002,
    g30869,g1003,g30870,g1004,g30871,g1005,g30713,g1006,g30714,g1007,g30715,
    g1009,g29635,g1010,g29636,g1008,g29637,g1090,g27206,g1091,g27207,g1089,
    g27208,g1137,g11536,g1138,g1139,g11537,g1140,g1141,g11538,g966,g967,g11518,
    g968,g969,g11519,g970,g971,g11520,g972,g973,g11521,g974,g975,g11522,g976,
    g977,g13423,g978,g986,g19024,g992,g27200,g995,g27201,g984,g27202,g983,
    g27203,g982,g27204,g981,g27205,g991,g19028,g990,g19027,g989,g19026,g988,
    g19025,g987,g25141,g985,g27199,g1029,g11524,g1036,g1037,g11525,g1038,g1039,
    g11526,g1040,g1044,g11527,g1051,g1052,g11528,g1053,g1054,g11529,g1055,
    g1059,g11530,g1066,g1067,g11531,g1068,g1069,g11532,g1070,g1074,g11533,
    g1081,g1082,g11534,g1083,g1084,g11535,g1011,g1012,g13424,g1018,g1024,g1231,
    g13435,g1237,g1236,g1240,g23198,g1243,g20560,g1196,g20561,g1199,g16469,
    g1209,g1210,g1250,g11539,g1255,g1256,g11542,g1257,g1258,g11543,g1259,g1260,
    g11544,g1251,g1252,g11540,g1253,g1254,g11541,g1176,g1161,g13425,g1168,
    g1172,g1173,g24333,g1174,g24334,g1175,g24335,g1142,g25150,g1145,g25142,
    g1148,g25143,g1164,g25147,g1165,g25148,g1166,g25149,g1167,g24330,g1171,
    g24331,g1151,g24332,g1152,g25144,g1155,g25145,g1158,g25146,g1214,g16470,
    g1221,g1228,g1229,g19033,g1230,g1234,g27217,g1235,g19034,g1186,g1244,
    g19035,g1245,g1262,g28245,g1263,g28246,g1261,g28247,g1265,g28248,g1266,
    g28249,g1264,g28250,g1268,g28251,g1269,g28252,g1267,g28253,g1271,g28254,
    g1272,g28255,g1270,g28256,g1273,g25994,g1276,g25995,g1279,g25996,g1282,
    g25997,g1285,g25998,g1288,g25999,g1300,g29143,g1303,g29144,g1306,g29145,
    g1291,g29140,g1294,g29141,g1297,g29142,g1177,g27209,g1180,g27210,g1183,
    g27211,g1192,g8293,g1193,g24336,g1194,g19029,g1195,g19030,g1200,g19031,
    g1201,g19032,g1202,g27216,g1203,g27215,g1204,g27214,g1205,g27213,g1206,
    g27212,g1211,g1215,g13426,g1216,g13427,g1217,g13428,g1218,g13429,g1219,
    g13430,g1220,g13431,g1222,g13432,g1223,g13433,g1224,g25993,g1227,g13434,
    g1309,g13436,g1312,g1315,g1316,g20562,g1345,g21944,g1326,g23199,g1319,
    g24337,g1339,g25151,g1332,g26000,g1346,g26708,g1358,g27218,g1352,g27698,
    g1365,g28257,g1372,g28682,g1378,g29146,g1385,g23200,g1386,g23201,g1384,
    g23202,g1388,g23203,g1389,g23204,g1387,g23205,g1391,g23206,g1392,g23207,
    g1390,g23208,g1394,g23209,g1395,g23210,g1393,g23211,g1397,g23212,g1398,
    g23213,g1396,g23214,g1400,g23215,g1401,g23216,g1399,g23217,g1403,g23218,
    g1404,g23219,g1402,g23220,g1406,g23221,g1407,g23222,g1405,g23223,g1409,
    g23224,g1410,g23225,g1408,g23226,g1412,g23227,g1413,g23228,g1411,g23229,
    g1415,g23230,g1416,g23231,g1414,g23232,g1418,g23233,g1419,g23234,g1417,
    g23235,g1421,g26709,g1422,g26710,g1420,g26711,g1424,g24338,g1425,g24339,
    g1423,g24340,g1520,g13437,g1517,g1547,g1512,g24341,g1513,g24342,g1511,
    g24343,g1515,g24344,g1516,g24345,g1514,g24346,g1524,g24347,g1525,g24348,
    g1523,g24349,g1527,g24350,g1528,g24351,g1526,g24352,g1530,g24353,g1531,
    g24354,g1529,g24355,g1533,g24356,g1534,g24357,g1532,g24358,g1536,g24359,
    g1537,g24360,g1535,g24361,g1539,g24362,g1540,g24363,g1538,g24364,g1542,
    g24365,g1543,g24366,g1541,g24367,g1545,g24368,g1546,g24369,g1544,g24370,
    g1551,g26713,g1552,g26714,g1550,g26715,g1554,g26716,g1555,g26717,g1553,
    g26718,g1557,g26719,g1558,g26720,g1556,g26721,g1560,g26722,g1561,g26723,
    g1559,g26724,g1567,g30536,g1570,g30537,g1573,g30538,g1612,g30878,g1615,
    g30879,g1618,g30880,g1576,g30872,g1579,g30873,g1582,g30874,g1621,g30881,
    g1624,g30882,g1627,g30883,g1585,g30539,g1588,g30540,g1591,g30541,g1630,
    g30545,g1633,g30546,g1636,g30547,g1594,g30542,g1597,g30543,g1600,g30544,
    g1639,g30548,g1642,g30549,g1645,g30550,g1603,g30875,g1606,g30876,g1609,
    g30877,g1648,g30884,g1651,g30885,g1654,g30886,g1466,g26001,g1462,g26712,
    g1457,g27219,g1453,g27699,g1448,g28258,g1444,g28683,g1439,g29147,g1435,
    g29427,g1430,g29641,g1426,g29802,g1562,g20563,g1564,g1563,g1657,g13438,
    g1786,g1782,g1690,g11550,g1735,g28259,g1724,g28260,g1727,g28261,g1750,
    g28262,g1739,g28263,g1742,g28264,g1765,g28265,g1754,g28266,g1757,g28267,
    g1779,g28268,g1769,g28269,g1772,g28270,g1789,g29434,g1792,g29435,g1795,
    g29436,g1798,g29645,g1801,g29646,g1804,g29647,g1808,g29437,g1809,g29438,
    g1807,g29439,g1810,g27700,g1813,g27701,g1816,g27702,g1819,g27703,g1822,
    g27704,g1825,g27705,g1829,g28684,g1830,g28685,g1828,g28686,g1693,g29803,
    g1694,g29804,g1695,g29805,g1696,g30887,g1697,g30888,g1698,g30889,g1699,
    g30716,g1700,g30717,g1701,g30718,g1703,g29642,g1704,g29643,g1702,g29644,
    g1784,g27221,g1785,g27222,g1783,g27223,g1831,g11563,g1832,g1833,g11564,
    g1834,g1835,g11565,g1660,g1661,g11545,g1662,g1663,g11546,g1664,g1665,
    g11547,g1666,g1667,g11548,g1668,g1669,g11549,g1670,g1671,g13439,g1672,
    g1680,g19036,g1686,g29428,g1689,g29429,g1678,g29430,g1677,g29431,g1676,
    g29432,g1675,g29433,g1685,g19040,g1684,g19039,g1683,g19038,g1682,g19037,
    g1681,g25152,g1679,g27220,g1723,g11551,g1730,g1731,g11552,g1732,g1733,
    g11553,g1734,g1738,g11554,g1745,g1746,g11555,g1747,g1748,g11556,g1749,
    g1753,g11557,g1760,g1761,g11558,g1762,g1763,g11559,g1764,g1768,g11560,
    g1775,g1776,g11561,g1777,g1778,g11562,g1705,g1706,g13440,g1712,g1718,g1925,
    g13451,g1931,g1930,g1934,g23236,g1937,g20564,g1890,g20565,g1893,g16471,
    g1903,g1904,g1944,g11566,g1949,g1950,g11569,g1951,g1952,g11570,g1953,g1954,
    g11571,g1945,g1946,g11567,g1947,g1948,g11568,g1870,g1855,g13441,g1862,
    g1866,g1867,g24374,g1868,g24375,g1869,g24376,g1836,g25161,g1839,g25153,
    g1842,g25154,g1858,g25158,g1859,g25159,g1860,g25160,g1861,g24371,g1865,
    g24372,g1845,g24373,g1846,g25155,g1849,g25156,g1852,g25157,g1908,g16472,
    g1915,g1922,g1923,g19045,g1924,g1928,g29445,g1929,g19046,g1880,g1938,
    g19047,g1939,g1956,g28271,g1957,g28272,g1955,g28273,g1959,g28274,g1960,
    g28275,g1958,g28276,g1962,g28277,g1963,g28278,g1961,g28279,g1965,g28280,
    g1966,g28281,g1964,g28282,g1967,g26003,g1970,g26004,g1973,g26005,g1976,
    g26006,g1979,g26007,g1982,g26008,g1994,g29151,g1997,g29152,g2000,g29153,
    g1985,g29148,g1988,g29149,g1991,g29150,g1871,g27224,g1874,g27225,g1877,
    g27226,g1886,g8302,g1887,g24377,g1888,g19041,g1889,g19042,g1894,g19043,
    g1895,g19044,g1896,g29444,g1897,g29443,g1898,g29442,g1899,g29441,g1900,
    g29440,g1905,g1909,g13442,g1910,g13443,g1911,g13444,g1912,g13445,g1913,
    g13446,g1914,g13447,g1916,g13448,g1917,g13449,g1918,g26002,g1921,g13450,
    g2003,g13452,g2006,g2009,g2010,g20566,g2039,g21945,g2020,g23237,g2013,
    g24378,g2033,g25162,g2026,g26009,g2040,g26725,g2052,g27227,g2046,g27706,
    g2059,g28283,g2066,g28687,g2072,g29154,g2079,g23238,g2080,g23239,g2078,
    g23240,g2082,g23241,g2083,g23242,g2081,g23243,g2085,g23244,g2086,g23245,
    g2084,g23246,g2088,g23247,g2089,g23248,g2087,g23249,g2091,g23250,g2092,
    g23251,g2090,g23252,g2094,g23253,g2095,g23254,g2093,g23255,g2097,g23256,
    g2098,g23257,g2096,g23258,g2100,g23259,g2101,g23260,g2099,g23261,g2103,
    g23262,g2104,g23263,g2102,g23264,g2106,g23265,g2107,g23266,g2105,g23267,
    g2109,g23268,g2110,g23269,g2108,g23270,g2112,g23271,g2113,g23272,g2111,
    g23273,g2115,g26726,g2116,g26727,g2114,g26728,g2118,g24379,g2119,g24380,
    g2117,g24381,g2214,g13453,g2211,g2241,g2206,g24382,g2207,g24383,g2205,
    g24384,g2209,g24385,g2210,g24386,g2208,g24387,g2218,g24388,g2219,g24389,
    g2217,g24390,g2221,g24391,g2222,g24392,g2220,g24393,g2224,g24394,g2225,
    g24395,g2223,g24396,g2227,g24397,g2228,g24398,g2226,g24399,g2230,g24400,
    g2231,g24401,g2229,g24402,g2233,g24403,g2234,g24404,g2232,g24405,g2236,
    g24406,g2237,g24407,g2235,g24408,g2239,g24409,g2240,g24410,g2238,g24411,
    g2245,g26730,g2246,g26731,g2244,g26732,g2248,g26733,g2249,g26734,g2247,
    g26735,g2251,g26736,g2252,g26737,g2250,g26738,g2254,g26739,g2255,g26740,
    g2253,g26741,g2261,g30551,g2264,g30552,g2267,g30553,g2306,g30896,g2309,
    g30897,g2312,g30898,g2270,g30890,g2273,g30891,g2276,g30892,g2315,g30899,
    g2318,g30900,g2321,g30901,g2279,g30554,g2282,g30555,g2285,g30556,g2324,
    g30560,g2327,g30561,g2330,g30562,g2288,g30557,g2291,g30558,g2294,g30559,
    g2333,g30563,g2336,g30564,g2339,g30565,g2297,g30893,g2300,g30894,g2303,
    g30895,g2342,g30902,g2345,g30903,g2348,g30904,g2160,g26010,g2156,g26729,
    g2151,g27228,g2147,g27707,g2142,g28284,g2138,g28688,g2133,g29155,g2129,
    g29446,g2124,g29648,g2120,g29806,g2256,g20567,g2258,g2257,g2351,g13454,
    g2480,g2476,g2384,g11577,g2429,g28285,g2418,g28286,g2421,g28287,g2444,
    g28288,g2433,g28289,g2436,g28290,g2459,g28291,g2448,g28292,g2451,g28293,
    g2473,g28294,g2463,g28295,g2466,g28296,g2483,g29447,g2486,g29448,g2489,
    g29449,g2492,g29652,g2495,g29653,g2498,g29654,g2502,g29450,g2503,g29451,
    g2501,g29452,g2504,g27708,g2507,g27709,g2510,g27710,g2513,g27711,g2516,
    g27712,g2519,g27713,g2523,g28689,g2524,g28690,g2522,g28691,g2387,g29807,
    g2388,g29808,g2389,g29809,g2390,g30905,g2391,g30906,g2392,g30907,g2393,
    g30719,g2394,g30720,g2395,g30721,g2397,g29649,g2398,g29650,g2396,g29651,
    g2478,g27230,g2479,g27231,g2477,g27232,g2525,g11590,g2526,g2527,g11591,
    g2528,g2529,g11592,g2354,g2355,g11572,g2356,g2357,g11573,g2358,g2359,
    g11574,g2360,g2361,g11575,g2362,g2363,g11576,g2364,g2365,g13455,g2366,
    g2374,g19048,g2380,g30314,g2383,g30315,g2372,g30316,g2371,g30317,g2370,
    g30318,g2369,g30319,g2379,g19052,g2378,g19051,g2377,g19050,g2376,g19049,
    g2375,g25163,g2373,g27229,g2417,g11578,g2424,g2425,g11579,g2426,g2427,
    g11580,g2428,g2432,g11581,g2439,g2440,g11582,g2441,g2442,g11583,g2443,
    g2447,g11584,g2454,g2455,g11585,g2456,g2457,g11586,g2458,g2462,g11587,
    g2469,g2470,g11588,g2471,g2472,g11589,g2399,g2400,g13456,g2406,g2412,g2619,
    g13467,g2625,g2624,g2628,g23274,g2631,g20568,g2584,g20569,g2587,g16473,
    g2597,g2598,g2638,g11593,g2643,g2644,g11596,g2645,g2646,g11597,g2647,g2648,
    g11598,g2639,g2640,g11594,g2641,g2642,g11595,g2564,g2549,g13457,g2556,
    g2560,g2561,g24415,g2562,g24416,g2563,g24417,g2530,g25172,g2533,g25164,
    g2536,g25165,g2552,g25169,g2553,g25170,g2554,g25171,g2555,g24412,g2559,
    g24413,g2539,g24414,g2540,g25166,g2543,g25167,g2546,g25168,g2602,g16474,
    g2609,g2616,g2617,g19057,g2618,g2622,g30325,g2623,g19058,g2574,g2632,
    g19059,g2633,g2650,g28297,g2651,g28298,g2649,g28299,g2653,g28300,g2654,
    g28301,g2652,g28302,g2656,g28303,g2657,g28304,g2655,g28305,g2659,g28306,
    g2660,g28307,g2658,g28308,g2661,g26012,g2664,g26013,g2667,g26014,g2670,
    g26015,g2673,g26016,g2676,g26017,g2688,g29159,g2691,g29160,g2694,g29161,
    g2679,g29156,g2682,g29157,g2685,g29158,g2565,g27233,g2568,g27234,g2571,
    g27235,g2580,g8311,g2581,g24418,g2582,g19053,g2583,g19054,g2588,g19055,
    g2589,g19056,g2590,g30324,g2591,g30323,g2592,g30322,g2593,g30321,g2594,
    g30320,g2599,g2603,g13458,g2604,g13459,g2605,g13460,g2606,g13461,g2607,
    g13462,g2608,g13463,g2610,g13464,g2611,g13465,g2612,g26011,g2615,g13466,
    g2697,g13468,g2700,g2703,g2704,g20570,g2733,g21946,g2714,g23275,g2707,
    g24419,g2727,g25173,g2720,g26018,g2734,g26742,g2746,g27236,g2740,g27714,
    g2753,g28309,g2760,g28692,g2766,g29162,g2773,g23276,g2774,g23277,g2772,
    g23278,g2776,g23279,g2777,g23280,g2775,g23281,g2779,g23282,g2780,g23283,
    g2778,g23284,g2782,g23285,g2783,g23286,g2781,g23287,g2785,g23288,g2786,
    g23289,g2784,g23290,g2788,g23291,g2789,g23292,g2787,g23293,g2791,g23294,
    g2792,g23295,g2790,g23296,g2794,g23297,g2795,g23298,g2793,g23299,g2797,
    g23300,g2798,g23301,g2796,g23302,g2800,g23303,g2801,g23304,g2799,g23305,
    g2803,g23306,g2804,g23307,g2802,g23308,g2806,g23309,g2807,g23310,g2805,
    g23311,g2809,g26743,g2810,g26744,g2808,g26745,g2812,g24420,g2813,g24421,
    g2811,g24422,g3054,g23317,g3079,g23318,g3080,g21965,g3043,g29453,g3044,
    g29454,g3045,g29455,g3046,g29456,g3047,g29457,g3048,g29458,g3049,g29459,
    g3050,g29460,g3051,g29655,g3052,g29972,g3053,g29973,g3055,g29974,g3056,
    g29975,g3057,g29976,g3058,g29977,g3059,g29978,g3060,g29979,g3061,g30119,
    g3062,g30908,g3063,g30909,g3064,g30910,g3065,g30911,g3066,g30912,g3067,
    g30913,g3068,g30914,g3069,g30915,g3070,g30940,g3071,g30980,g3072,g30981,
    g3073,g30982,g3074,g30983,g3075,g30984,g3076,g30985,g3077,g30986,g3078,
    g30987,g2997,g30989,g2993,g26748,g2998,g27238,g3006,g25177,g3002,g26021,
    g3013,g26750,g3010,g27239,g3024,g27716,g3018,g24425,g3028,g25176,g3036,
    g26022,g3032,g26749,g3040,g16497,g2986,g2987,g16495,g48,g20595,g45,g20596,
    g42,g20597,g39,g20598,g27,g20599,g30,g20600,g33,g20601,g36,g20602,g3083,
    g20603,g26,g20604,g2992,g21966,g23,g20605,g20,g20606,g17,g20607,g11,g20608,
    g14,g20589,g5,g20590,g8,g20591,g2,g20592,g2990,g20593,g2991,g21964,g1,
    g20594,II13089,g562,II13092,g1248,II13095,g1942,II13098,g2636,II13101,
    g3235,II13104,g3236,II13107,g3237,II13110,g3238,II13113,g3239,II13116,
    g3240,II13119,g3241,II13122,g3242,II13125,g3243,II13128,g3244,II13131,
    g3245,II13134,g3246,II13137,g3247,II13140,g3248,II13143,g3249,II13146,
    g3250,II13149,g3251,II13152,g3252,II13155,g3253,II13158,g3254,II13161,
    g3304,g3305,II13165,g3306,g3337,II13169,g3338,g3365,II13173,g3366,II13176,
    g3398,II13179,g3410,II13182,g3460,g3461,II13186,g3462,g3493,II13190,g3494,
    g3521,II13194,g3522,II13197,g3554,II13200,g3566,II13203,g3616,g3617,
    II13207,g3618,g3649,II13211,g3650,g3677,II13215,g3678,II13218,g3710,
    II13221,g3722,II13224,g3772,g3773,II13228,g3774,g3805,II13232,g3806,g3833,
    II13236,g3834,II13239,g3866,II13242,g3878,g3897,II13246,g3900,g3919,g3922,
    g3925,g3928,g3931,g3934,g3937,g3940,g3941,g3942,g3945,g3948,g3951,g3954,
    g3957,g3960,g3963,g3966,g3969,g3972,g3975,g3978,g3981,g3984,g3987,g3990,
    II13275,g3994,g3995,g3996,g3997,g3998,g3999,g4000,g4003,g4006,g4009,g4012,
    g4015,g4016,g4017,g4020,g4023,g4026,g4029,g4032,g4035,g4038,g4041,g4044,
    g4047,g4048,g4049,g4052,g4055,g4058,g4061,g4064,g4067,g4070,g4073,g4076,
    g4079,g4082,g4085,II13316,g4089,II13320,g4091,g4092,g4093,g4094,g4095,
    g4098,g4101,g4104,g4107,g4110,g4111,g4112,g4115,g4118,g4121,g4124,g4127,
    g4130,g4133,g4136,g4139,g4142,g4143,g4144,g4147,g4150,g4153,g4156,g4159,
    g4162,g4165,g4168,g4171,g4174,g4175,g4176,g4179,g4182,g4185,g4188,g4191,
    g4194,g4197,II13366,g4201,g4202,g4203,g4204,g4205,g4208,g4211,g4214,g4217,
    g4220,g4221,g4224,g4225,g4228,g4231,g4234,g4237,g4240,g4243,g4246,g4249,
    g4250,g4251,g4254,g4257,g4260,g4263,g4266,g4269,g4272,g4275,g4278,g4281,
    g4282,g4283,g4286,g4289,g4292,g4295,g4298,g4301,g4304,g4307,g4310,g4313,
    g4314,g4315,g4318,II13417,g4322,II13421,g4324,g4325,g4326,g4329,g4332,
    g4335,II13430,g4338,II13433,g4339,g4340,g4343,g4346,g4347,g4348,g4351,
    g4354,g4357,g4360,g4363,g4366,g4369,g4372,g4375,g4376,g4379,g4380,g4383,
    g4386,g4389,g4392,g4395,g4398,g4401,g4404,g4405,g4406,g4409,g4412,g4415,
    g4418,g4421,g4424,g4427,g4430,g4433,g4436,g4437,g4438,g4441,g4444,g4447,
    II13478,g4451,g4452,g4453,g4456,g4465,g4468,g4471,g4474,g4475,g4476,g4479,
    g4480,g4483,g4486,g4489,g4492,g4495,g4498,g4501,g4504,II13501,g4507,
    II13504,g4508,g4509,g4512,g4515,g4516,g4517,g4520,g4523,g4526,g4529,g4532,
    g4535,g4538,g4541,g4544,g4545,g4548,g4549,g4552,g4555,g4558,g4561,g4564,
    g4567,g4570,g4573,g4574,g4575,g4578,g4581,g4584,g4587,II13538,g4591,g4592,
    g4595,g4598,g4601,g4602,g4603,g4606,g4609,g4610,g4611,g4614,g4617,g4620,
    g4623,g4626,g4629,g4632,g4641,g4644,g4647,g4650,g4651,g4652,g4655,g4656,
    g4659,g4662,g4665,g4668,g4671,g4674,g4677,g4680,II13575,g4683,II13578,
    g4684,g4685,g4688,g4691,g4692,g4693,g4696,g4699,g4702,g4705,g4708,g4711,
    g4714,g4717,g4720,g4721,g4724,g4725,g4728,g4731,g4734,II13601,g4735,
    II13604,g4736,g4737,g4740,g4743,g4746,g4749,g4752,g4753,g4754,g4757,g4760,
    g4763,g4766,g4769,g4772,g4775,g4778,g4779,g4780,g4783,g4786,g4787,g4788,
    g4791,g4794,g4797,g4800,g4803,g4806,g4809,g4818,g4821,g4824,g4827,g4828,
    g4829,g4832,g4833,g4836,g4839,g4842,g4845,g4848,g4851,g4854,g4857,II13652,
    g4860,II13655,g4861,g4862,g4865,g4868,g4869,g4870,g4873,g4876,g4879,g4882,
    g4885,g4888,g4891,g4894,g4897,g4898,g4899,g4902,g4905,g4908,II13677,g4911,
    II13680,g4912,g4913,g4916,g4919,g4922,g4925,g4928,g4929,g4930,g4933,g4936,
    g4939,g4942,g4945,g4948,g4951,g4954,g4955,g4956,g4959,g4962,g4963,g4964,
    g4967,g4970,g4973,g4976,g4979,g4982,g4985,g4994,g4997,g5000,g5003,g5004,
    g5005,g5008,g5009,g5012,g5015,g5018,g5021,g5024,g5027,g5030,g5033,g5034,
    g5035,g5038,g5041,g5044,g5047,g5050,g5053,g5056,g5057,g5058,g5061,g5064,
    g5067,II13742,g5070,II13745,g5071,g5072,g5075,g5078,g5081,g5084,g5087,
    g5088,g5089,g5092,g5095,g5098,g5101,g5104,g5107,g5110,g5113,g5114,g5115,
    g5118,g5121,g5122,g5123,g5126,g5129,g5132,g5135,g5138,II13775,g5141,g5142,
    g5145,g5148,g5149,g5150,g5153,g5156,g5159,g5162,g5163,g5164,g5167,g5170,
    g5173,g5176,g5179,g5182,g5185,g5186,g5187,g5190,g5193,g5196,II13801,g5199,
    II13804,g5200,g5201,g5204,g5207,g5210,g5213,g5216,g5217,g5218,g5221,g5224,
    g5227,g5230,g5233,II13820,g5234,g5235,g5238,g5241,g5242,g5243,g5246,g5249,
    g5252,g5255,g5256,g5257,g5260,g5263,g5266,g5269,g5272,g5275,g5278,g5279,
    g5280,g5283,g5286,g5289,g5292,g5293,g5296,II13849,g5297,g5298,g5301,g5304,
    g5305,g5306,g5309,g5312,g5315,g5318,g5319,g5320,g5323,g5326,g5327,g5330,
    g5333,II13868,g5334,g5335,g5338,g5341,g5342,g5343,g5346,g5349,g5352,g5355,
    g5358,g5361,g5362,g5363,g5366,g5369,g5372,g5375,g5378,g5379,g5382,g5385,
    II13892,g5389,II13896,g5390,g5391,g5394,II13901,g5395,II13904,g5396,
    II13907,g5397,II13910,g5398,II13913,g5399,II13916,g5400,II13919,g5401,
    II13922,g5402,II13925,g5403,II13928,g5404,II13931,g5405,II13934,g5406,
    II13937,g5407,II13940,g5408,II13943,g5409,g5410,II13947,g5411,II13950,
    g5412,II13953,g5413,II13956,g5414,II13959,g5415,II13962,g5416,II13965,
    g5417,II13968,g5418,II13971,g5419,II13974,g5420,II13977,g5421,II13980,
    g5422,g5423,II13984,g5424,II13987,g5425,II13990,g5426,II13993,g5427,g5428,
    g5431,g5434,II13999,II14002,g5438,g5469,II14006,II14009,g5473,g5504,g5507,
    II14014,g5508,II14017,II14020,g5512,g5543,g5546,g5547,g5548,II14027,
    II14030,g5550,g5551,II14034,g5552,II14037,II14040,g5556,g5587,g5590,g5591,
    g5592,g5593,g5594,II14049,II14052,g5596,g5597,II14056,g5598,g5601,g5604,
    g5605,g5606,g5609,g5610,g5611,II14066,II14069,g5613,g5614,II14073,g5615,
    g5618,g5621,g5622,g5623,g5626,g5627,g5628,II14083,g5631,g5634,g5635,g5636,
    II14091,II14094,g5638,g5639,g5640,g5641,g5642,g5645,g5646,g5647,II14104,
    g5651,g5654,g5655,g5656,II14113,g5659,g5662,g5663,g5664,g5665,g5666,g5667,
    g5668,g5675,g5679,g5680,g5683,g5684,g5685,II14134,g5689,g5692,g5693,g5694,
    II14143,g5697,g5700,II14149,g5701,g5702,g5703,g5704,g5705,g5706,g5707,
    g5708,g5712,II14163,g5713,g5714,g5715,g5716,g5717,g5718,g5719,g5720,g5727,
    g5731,g5732,g5735,g5736,g5737,II14182,g5741,g5744,g5745,g5746,II14191,
    II14195,g5749,g5750,g5751,g5752,g5753,g5754,g5755,g5756,g5759,g5760,g5761,
    g5762,g5763,g5764,g5765,g5766,g5770,II14219,g5771,g5772,g5773,g5774,g5775,
    g5776,g5777,g5778,g5785,g5789,g5790,g5793,g5794,g5795,II14238,II14243,
    g5799,II14246,g5800,II14249,g5801,g5802,g5803,g5804,g5805,g5806,g5808,
    g5809,g5810,g5811,g5812,g5813,g5814,g5815,g5818,g5819,g5820,g5821,g5822,
    g5823,g5824,g5825,g5829,II14280,g5830,g5831,g5832,g5833,g5834,g5835,g5836,
    g5837,g5844,g5848,II14295,g5849,II14298,g5850,g5851,g5852,g5853,g5854,
    g5855,II14306,g5856,g5857,g5858,g5859,g5860,g5861,g5862,g5864,g5865,g5866,
    g5867,g5868,g5869,g5870,g5871,g5874,g5875,g5876,g5877,g5878,g5879,g5880,
    g5881,g5885,II14338,g5886,g5887,g5888,II14343,g5889,g5890,g5893,g5894,
    g5895,g5896,g5897,g5898,g5899,g5900,g5901,g5902,II14357,g5903,g5904,g5905,
    g5906,g5907,g5908,g5909,g5911,g5912,g5913,g5914,g5915,g5916,g5917,g5918,
    g5921,II14378,g5922,II14381,g5923,II14384,g5924,g5925,g5926,g5927,g5928,
    g5929,g5932,g5933,g5934,g5935,g5936,g5937,g5938,g5939,g5940,g5941,II14402,
    g5942,g5943,g5944,g5945,g5946,g5947,g5948,g5950,II14413,g5951,II14416,
    g5952,g5953,g5954,g5955,g5956,g5957,II14424,g5958,g5959,g5960,g5961,g5962,
    g5963,g5966,g5967,g5968,g5969,g5970,g5971,g5972,g5973,g5974,g5975,II14442,
    g5976,g5977,II14446,g5978,II14449,g5979,g5980,g5981,g5982,g5983,g5984,
    g5985,g5986,II14459,g5987,g5988,g5989,g5990,g5991,g5992,g5995,g5996,g5997,
    g5998,g5999,II14472,g6000,II14475,g6014,II14478,g6015,g6016,g6017,g6018,
    g6019,g6020,g6021,g6022,g6023,II14489,g6024,g6025,g6026,g6027,g6028,
    II14496,g6029,II14499,g6030,II14502,g6031,g6032,g6033,g6034,g6035,g6036,
    g6037,g6038,g6039,II14513,g6040,II14516,g6041,II14519,g6042,g6043,g6044,
    g6045,II14525,g6046,g6047,II14529,g6048,II14532,g6051,II14535,g6052,
    II14538,g6053,II14541,g6054,II14544,g6055,II14547,g6056,II14550,g6057,
    II14553,g6058,II14556,g6059,II14559,g6060,II14562,g6061,II14565,g6062,
    II14568,g6063,II14571,g6064,II14574,g6065,II14577,g6066,II14580,g6067,
    g6068,II14584,g6079,II14587,g6080,II14590,g6081,II14593,g6082,II14596,
    g6083,II14599,g6084,II14602,g6085,II14605,g6086,g6087,II14609,g6098,
    II14612,g6099,II14615,g6100,II14618,g6101,II14621,g6102,II14624,g6103,
    g6104,II14628,g6115,II14631,g6116,II14634,g6117,II14637,g6118,g6119,
    II14641,g6130,II14644,g6131,II14647,g6134,II14650,g6135,g6136,II14654,
    g6139,g6140,g6141,g6142,II14660,g6145,g6146,g6149,II14665,g6153,II14668,
    g6156,g6157,g6161,g6162,g6163,II14675,g6166,g6167,g6170,g6173,g6177,g6180,
    g6183,g6184,g6188,g6189,g6190,II14688,g6193,g6194,g6197,g6200,g6201,g6204,
    g6205,g6209,g6212,g6215,g6216,g6220,g6221,g6222,II14704,g6226,g6227,
    II14709,g6230,II14712,II14715,g6232,g6281,g6284,g6288,g6289,g6290,g6293,
    g6294,g6298,g6301,g6304,g6305,g6309,g6310,II14731,II14734,g6314,g6363,
    g6367,II14739,II14742,g6369,g6418,g6421,g6425,g6426,g6427,g6430,g6431,
    g6435,g6438,g6441,II14755,g6443,g6444,II14760,II14763,g6448,II14766,
    II14769,g6486,g6512,g6513,g6517,II14775,II14778,g6519,g6568,g6572,II14783,
    II14786,g6574,g6623,g6626,g6630,g6631,g6632,g6635,g6636,g6637,g6638,g6641,
    II14799,II14802,g6643,g6672,g6675,g6676,II14808,II14811,g6678,g6707,g6711,
    II14816,II14819,g6713,II14822,II14825,g6751,g6776,g6777,g6781,II14831,
    II14834,g6783,g6832,g6836,II14839,II14842,g6838,g6887,g6890,g6894,II14848,
    g6896,g6897,g6898,g6901,g6905,g6908,II14857,II14860,g6912,g6942,g6943,
    II14865,II14868,g6945,g6974,g6977,g6978,II14874,II14877,g6980,g7009,g7013,
    II14882,II14885,g7015,II14888,II14891,g7053,g7078,g7079,g7083,II14897,
    II14900,g7085,g7134,g7138,g7139,g7140,g7141,g7142,g7143,g7146,g7149,g7152,
    g7153,g7156,g7157,g7158,II14917,II14920,g7162,g7192,g7193,II14925,II14928,
    g7195,g7224,g7227,g7228,II14934,II14937,g7230,g7259,g7263,II14942,II14945,
    g7265,II14948,II14951,g7303,g7328,g7329,g7333,II14957,g7335,g7336,g7337,
    g7338,g7342,g7345,g7346,g7347,g7348,g7349,g7352,g7353,g7354,II14973,
    II14976,g7358,g7388,g7389,II14981,II14984,g7391,g7420,g7423,g7424,II14990,
    II14993,g7426,g7455,g7459,g7460,g7461,g7462,g7465,g7466,g7471,g7475,g7476,
    g7477,g7478,g7479,g7482,g7483,g7484,II15012,II15015,g7488,g7518,II15019,
    g7520,g7521,g7522,g7527,g7529,g7530,g7531,g7532,g7533,g7534,g7535,g7538,
    g7539,g7540,g7541,g7542,g7545,g7548,g7549,g7553,g7554,g7555,g7556,g7557,
    g7558,g7559,g7560,g7561,g7562,g7566,g7570,g7573,g7574,g7576,g7577,g7578,
    g7579,g7580,g7581,g7582,g7583,g7587,g7590,g7591,g7592,g7593,g7594,g7595,
    g7600,g7603,g7604,g7605,g7606,g7607,g7610,g7613,g7614,g7615,g7616,g7619,
    g7622,g7623,g7626,g7629,g7632,g7635,g7638,g7639,g7642,g7643,g7646,g7649,
    g7652,g7655,g7658,g7661,g7664,g7667,g7670,g7673,g7676,g7679,g7682,g7685,
    g7688,g7691,g7694,g7697,g7700,g7703,g7706,g7709,g7712,g7715,g7718,g7721,
    g7724,g7727,g7730,g7733,g7736,g7739,g7742,g7745,g7748,g7751,g7754,g7757,
    g7760,g7763,g7766,g7769,g7772,g7776,g7779,g7782,g7785,g7788,g7792,g7796,
    g7799,g7802,g7806,g7809,g7812,g7815,g7819,g7822,g7823,g7826,g7827,g7830,
    g7833,g7834,g7837,g7838,g7841,g7842,g7845,g7848,g7849,g7852,g7856,g7857,
    g7858,g7861,g7862,g7865,g7868,g7869,g7872,g7877,g7878,g7879,g7880,g7888,
    g7891,g7892,g7897,g7898,g7899,g7900,II15222,g7901,g7906,II15226,g7910,
    II15230,g7911,g7912,g7915,g7916,g7919,g7924,g7925,g7926,g7927,g7928,
    II15256,g7936,g7949,g7950,g7953,II15262,g7957,g7958,II15267,g7962,II15271,
    g7963,g7964,g7967,g7971,g7972,g7973,g7974,g7975,II15288,g7976,g7989,g7990,
    g7993,g7996,g7999,g8000,g8001,g8004,II15299,g8008,g8009,II15304,g8013,
    II15308,g8014,g8015,g8018,II15313,g8022,II15317,g8024,g8025,g8026,g8027,
    g8028,g8029,II15326,II15329,g8031,g8044,g8045,g8053,g8056,g8059,g8062,
    g8065,g8068,g8071,g8074,g8075,g8076,g8079,II15345,g8083,g8084,II15350,
    g8088,II15354,g8089,g8090,g8093,II15359,g8097,g8098,g8099,g8100,g8101,
    g8102,g8103,II15369,II15372,g8107,g8120,g8123,g8126,g8129,g8132,g8135,
    g8138,g8141,g8144,g8147,g8150,g8153,g8156,g8159,g8160,g8161,g8164,II15392,
    g8168,g8169,g8172,II15398,g8176,g8177,g8178,g8179,g8180,g8181,g8182,g8183,
    g8191,g8194,g8197,g8200,g8203,g8206,g8209,g8212,g8215,g8218,g8221,g8224,
    g8227,g8230,g8233,g8236,g8239,g8242,g8245,g8246,II15429,g8250,II15433,
    g8252,g8253,g8254,g8255,g8256,g8257,II15442,II15445,II15448,II15451,
    II15454,II15457,II15460,II15463,II15466,II15469,II15472,II15475,II15478,
    II15481,II15484,II15487,II15490,II15493,g8276,g8277,g8278,II15499,g8285,
    g8286,g8287,II15505,g8294,g8295,g8296,II15511,g8303,g8304,g8305,II15517,
    g8312,g8313,g8317,II15523,g8321,II15526,g8324,II15532,g8330,II15535,g8333,
    II15538,g8336,II15543,g8341,II15546,g8344,II15549,g8347,II15553,g8351,
    II15556,g8354,II15559,g8357,II15562,g8360,II15565,g8363,II15568,g8366,
    II15571,g8369,II15574,g8372,II15577,g8375,II15580,g8378,II15584,g8382,
    II15590,g8388,II15593,g8391,II15599,g8397,II15602,g8400,II15605,g8403,
    II15610,g8408,II15613,g8411,II15616,g8414,II15620,g8418,II15623,g8421,
    II15626,g8424,II15629,g8427,II15636,g8434,II15642,g8440,II15645,g8443,
    II15651,g8449,II15654,g8452,II15657,g8455,II15662,g8460,II15671,g8469,
    II15677,g8475,II15680,g8478,II15696,g8494,g8514,g8530,g8568,II15771,g8569,
    II15779,g8575,II15784,g8578,II15787,g8579,g8580,g8587,g8594,II15794,g8602,
    g8605,II15800,g8614,II15803,g8617,II15806,g8620,II15810,g8622,II15815,
    g8627,II15818,g8630,II15822,g8632,II15827,g8637,II15830,g8640,II15833,
    g8643,II15836,g8646,II15839,g8649,II15843,g8651,II15847,g8655,II15850,
    g8658,II15853,g8659,II15856,g8662,II15859,g8665,II15863,g8667,II15866,
    g8670,II15869,g8673,II15873,g8677,II15876,g8678,II15879,g8681,II15882,
    g8684,II15887,g8689,II15890,g8690,II15893,g8693,II15896,g8696,II15899,
    g8699,II15902,g8700,II15909,g8707,II15912,g8708,II15915,g8711,II15918,
    g8714,II15922,g8718,II15925,g8719,II15932,g8726,II15935,g8745,II15938,
    g8748,II15942,g8752,II15946,g8756,II15949,g8757,II15955,g8763,II15958,
    g8766,II15961,g8769,II15964,g8770,II15967,g8771,II15971,g8775,II15975,
    g8779,II15978,g8780,II15983,g8785,II15986,g8788,II15989,g8791,II15992,
    g8792,II15995,g8793,II15998,g8794,II16002,g8798,II16006,g8802,II16009,
    g8805,II16012,g8808,II16015,g8809,II16018,g8810,II16021,g8811,II16024,
    g8812,II16027,g8813,II16031,g8817,II16034,g8820,II16037,g8821,g8822,
    II16041,g8823,II16044,g8824,II16047,g8825,II16050,g8826,II16053,g8827,
    II16056,g8828,II16059,g8829,II16062,g8832,II16065,g8835,II16068,g8836,
    II16071,g8839,II16074,g8840,II16079,g8843,II16082,g8844,II16085,g8845,
    g8846,II16089,g8847,II16092,g8850,II16095,g8851,II16098,g8852,II16101,
    g8853,II16104,g8856,II16107,g8859,II16110,g8860,II16114,g8862,II16117,
    g8863,II16120,g8866,II16123,g8867,II16128,g8870,II16131,g8871,II16134,
    g8872,g8873,II16138,g8874,II16141,g8877,II16144,g8878,II16147,g8879,
    II16150,g8882,II16153,g8885,II16156,g8888,II16159,g8891,II16163,g8893,
    II16166,g8894,II16169,g8897,II16172,g8898,II16176,g8900,II16179,g8901,
    II16182,g8904,II16185,g8905,II16190,g8908,II16193,g8909,II16196,g8910,
    g8911,II16200,g8912,II16203,g8915,II16206,g8918,II16209,g8921,II16212,
    g8924,II16215,g8925,II16218,g8928,II16221,g8931,II16225,g8933,II16228,
    g8934,II16231,g8937,II16234,g8938,II16238,g8940,II16241,g8941,II16244,
    g8944,II16247,g8945,II16252,g8948,II16255,g8949,II16258,g8952,II16261,
    g8955,II16264,g8958,II16267,g8961,II16270,g8964,II16273,g8965,II16276,
    g8968,II16279,g8971,II16283,g8973,II16286,g8974,II16289,g8977,II16292,
    g8978,II16296,g8980,g8983,II16300,g8984,II16303,g8987,II16306,g8990,
    II16309,g8993,II16312,g8996,II16315,g8997,II16318,g9000,II16321,g9003,
    II16325,g9005,II16328,g9006,II16332,g9010,II16335,g9013,II16338,g9016,
    II16341,g9019,II16344,g9022,II16347,g9025,g9027,II16354,g9035,II16357,
    g9038,II16360,g9041,II16363,g9044,g9050,II16372,g9058,g9067,g9084,II16432,
    g9128,II16438,g9134,II16444,g9140,II16450,g9146,II16453,g9149,g9150,
    II16457,g9159,g9160,g9161,II16462,g9170,II16465,g9173,g9174,II16469,g9183,
    II16472,g9184,g9187,II16476,g9196,II16479,g9199,II16482,g9202,g9203,
    II16486,g9212,II16489,g9215,g9216,II16493,g9225,g9226,g9227,g9228,II16499,
    g9229,g9232,II16504,g9242,II16507,g9245,g9248,II16511,g9257,II16514,g9260,
    II16517,g9263,g9264,II16521,g9273,II16524,g9276,g9277,g9286,g9287,g9288,
    g9289,II16532,g9290,g9293,II16538,g9303,II16541,g9306,II16544,g9309,g9310,
    II16549,g9320,II16552,g9323,g9326,II16556,g9335,II16559,g9338,II16562,
    g9341,g9342,II16566,g9351,II16569,g9354,g9355,g9356,II16578,g9368,II16581,
    g9371,g9374,II16587,g9384,II16590,g9387,II16593,g9390,g9391,II16598,g9401,
    II16601,g9404,g9407,II16605,g9416,II16608,g9419,II16611,g9422,g9423,g9424,
    g9425,g9426,g9427,II16624,g9443,II16627,g9446,II16630,g9449,II16633,g9450,
    g9453,II16641,g9465,II16644,g9468,g9471,II16650,g9481,II16653,g9484,
    II16656,g9487,g9488,II16661,g9498,II16664,g9501,g9504,g9505,g9506,g9507,
    II16677,g9524,g9527,II16681,g9528,II16684,g9531,g9569,II16694,g9585,
    II16697,g9588,II16700,g9591,II16703,g9592,g9595,II16711,g9607,II16714,
    g9610,g9613,II16720,g9623,II16723,g9626,II16726,g9629,II16741,g9640,
    II16744,g9641,II16747,g9644,g9649,II16759,g9666,g9669,II16763,g9670,
    II16766,g9673,g9711,II16776,g9727,II16779,g9730,II16782,g9733,II16785,
    g9734,g9737,II16793,g9749,II16796,g9752,g9755,g9756,g9757,g9758,II16811,
    g9767,II16814,g9770,II16832,g9786,II16835,g9787,II16838,g9790,g9795,
    II16850,g9812,g9815,II16854,g9816,II16857,g9819,g9857,II16867,g9873,
    II16870,g9876,II16873,g9879,II16876,g9880,g9884,g9885,g9886,II16897,g9895,
    II16900,g9898,II16915,g9913,II16918,g9916,II16936,g9932,II16939,g9933,
    II16942,g9936,g9941,II16954,g9958,g9961,II16958,g9962,II16961,g9965,
    II16972,g10004,g10015,II16984,g10016,II16987,g10017,II16990,g10018,II16993,
    g10021,II17009,g10049,II17012,g10052,II17027,g10067,II17030,g10070,II17048,
    g10086,II17051,g10087,II17054,g10090,II17066,g10096,g10099,II17070,g7528,
    g10100,II17081,g10109,g10124,II17097,g10125,II17100,g10126,II17103,g10127,
    II17106,g10130,II17122,g10158,II17125,g10161,II17140,g10176,II17143,g10179,
    II17159,g10189,II17184,g10214,g10229,II17200,g10230,II17203,g10231,II17206,
    g10232,II17209,g10235,II17225,g10263,II17228,g10266,II17235,g10273,II17238,
    g10276,II17278,g10316,g10331,II17294,g10332,II17297,g10333,II17300,g10334,
    II17303,g10337,II17311,g10357,II17363,g10409,II17370,g10416,II17373,g10419,
    g10424,g10481,II17433,g10482,g10486,g10500,II17483,g10542,II17486,g10545,
    g10549,g10560,g10574,II17527,g10601,g10606,g10617,g10631,II17557,g10646,
    g10653,g10664,g10683,g10694,g10714,g10730,g10735,g10749,g10754,g10765,
    g10766,g10767,g10772,g10773,II17627,g7575,g10779,g10783,II17632,g10787,
    g10788,II17637,g10792,II17641,g10796,II17645,g10800,II17649,g10804,II17653,
    g10808,g10809,II17658,g10813,II17662,g10817,II17666,g10821,II17670,g10825,
    II17673,g10826,g10829,II17677,g10830,II17681,g10834,II17685,g10838,II17689,
    g10842,II17692,g10843,g10846,g10847,g10848,II17698,g10849,II17701,g10850,
    II17705,g10854,II17709,g10858,II17712,g10859,II17715,g10862,g10865,g10866,
    g10867,II17721,g10868,II17724,g10869,II17727,g10870,II17730,g10871,II17734,
    g10875,II17737,g10876,II17740,g10877,II17743,g10880,II17746,g10883,g10886,
    II17750,g10887,II17753,g10888,II17756,g10889,II17759,g10890,II17762,g10891,
    II17765,g10892,II17768,g10895,II17771,g10898,II17774,g10901,g10904,g10905,
    g10906,II17780,g10907,II17783,g10908,II17786,g10909,II17789,g10910,II17792,
    g10911,II17795,g10912,II17798,g10915,II17801,g10918,II17804,g10921,II17807,
    g10924,g10927,g10928,g10929,II17813,g10930,II17816,g10931,II17819,g10932,
    II17822,g10933,II17825,g10934,II17828,g10935,II17831,g10936,II17834,g10937,
    II17837,g10940,II17840,g10943,II17843,g10946,II17846,g10949,II17849,g10952,
    g10961,g10962,II17854,g10963,II17857,g10966,II17860,g10967,II17863,g10968,
    II17866,g10969,II17869,g10972,II17872,g10973,II17875,g10974,II17878,g10977,
    II17881,g10980,II17884,g10983,g10986,g10987,II17889,g10988,II17892,g10991,
    II17895,g10994,II17898,g10995,II17901,g10996,II17904,g10999,II17907,g11002,
    II17910,g11003,II17913,g11004,II17916,g11007,II17919,g11008,II17922,g11011,
    II17925,g11014,II17928,g11017,g11020,g11021,II17933,g11022,II17936,g11025,
    II17939,g11028,II17942,g11031,II17945,g11032,II17948,g11035,II17951,g11036,
    II17954,g11039,II17957,g11042,II17960,g11045,II17963,g11048,II17966,g11051,
    II17969,g11054,II17972,g11055,II17975,g11056,II17978,g7795,g11059,II17981,
    g11063,II17984,g11066,g11069,g11078,II17989,g11079,II17992,g11082,II17995,
    g11085,II17998,g11088,II18001,g11091,II18004,g11092,II18007,g11095,II18010,
    g11098,II18013,g11101,II18016,g11102,II18019,g11105,II18022,g11108,II18025,
    g11111,II18028,g11114,II18031,g11117,II18034,g11120,II18037,g11123,II18040,
    g11126,II18043,g11129,II18046,g11132,II18049,g11135,II18052,g11138,II18055,
    g11141,II18058,g11144,II18061,g11145,II18064,g11148,II18067,g11151,II18070,
    g11154,II18073,g11157,II18076,g11160,II18079,g11163,II18082,g11166,II18085,
    g11169,II18088,g11170,II18091,g11173,II18094,g11176,II18097,g11179,II18100,
    g11182,II18103,g11185,g11190,II18121,g11199,II18124,g11202,II18127,g11205,
    II18130,g11208,II18133,g11209,II18136,g11210,II18139,g11213,II18142,g11216,
    II18145,g11219,II18148,g11222,II18151,g11225,II18154,g11228,II18157,g11231,
    II18160,g11234,II18163,g11237,II18166,g11240,II18169,g11243,II18172,g11246,
    II18175,g11249,II18178,g11252,II18181,g11255,II18184,g11256,II18187,g11259,
    II18211,g11265,II18214,g11268,II18217,g11271,II18220,g11274,II18223,g11277,
    II18226,g11278,II18229,g11281,II18232,g11284,II18235,g11287,II18238,g11290,
    II18241,g11291,II18244,g11294,II18247,g11297,II18250,g11300,II18253,g11303,
    II18256,g11306,II18259,g11309,II18262,g11312,II18265,g11315,II18268,g11318,
    II18271,g11321,II18274,g11324,II18277,g11327,g11332,II18295,g11341,II18298,
    g11344,II18302,g11348,II18305,g11351,II18308,g11354,II18311,g11355,II18314,
    g11358,II18317,g11361,II18320,g11364,II18323,g11367,II18326,g11370,II18329,
    g11373,II18332,g11376,II18335,g11379,II18338,g11382,II18341,g11385,II18344,
    g11386,II18347,g11389,II18350,g11392,II18353,g11395,II18356,g11398,II18359,
    g11401,II18362,g11404,II18365,g11407,II18375,g11411,II18378,g11414,II18381,
    g11417,II18386,g11422,II18389,g11425,II18392,g11428,II18396,g11432,II18399,
    g11435,II18402,g11438,II18405,g11441,II18408,g11444,II18411,g11447,II18414,
    g11450,II18417,g11453,II18420,g11456,II18423,g11459,II18426,g11462,II18429,
    g11465,II18432,g11468,II18435,g11471,II18438,g11472,II18441,g11475,II18444,
    g11478,g11481,g11490,II18449,II18452,II18455,II18458,II18461,II18464,
    II18467,II18470,II18473,II18476,II18479,II18482,II18485,II18488,II18491,
    II18494,II18497,II18500,II18503,II18506,II18509,II18512,II18515,II18518,
    II18521,II18524,II18527,II18530,II18533,II18536,II18539,II18542,II18545,
    II18548,II18551,II18554,II18557,II18560,II18563,II18566,II18569,II18572,
    II18575,II18578,II18581,II18584,II18587,II18590,II18593,II18596,II18599,
    II18602,II18605,II18608,II18611,II18614,II18617,II18620,II18623,II18626,
    II18629,II18632,II18635,II18638,II18641,II18644,II18647,II18650,II18653,
    II18656,II18659,II18662,II18665,II18668,II18671,II18674,II18677,II18680,
    II18683,II18686,II18689,II18692,II18695,II18698,II18701,II18704,II18707,
    II18710,II18713,II18716,II18719,II18722,II18725,II18728,II18731,II18734,
    II18737,II18740,II18743,II18746,II18749,II18752,II18755,II18758,II18761,
    II18764,II18767,II18770,II18773,g11599,II18777,g11603,II18780,g11606,
    II18784,g11608,II18787,g11611,II18791,g11613,II18794,g11616,g11620,g11623,
    II18810,g11628,II18813,g11629,II18817,g11633,II18820,g11636,II18824,g11638,
    II18827,g11641,g11642,II18835,g11651,II18838,g11652,II18842,g11656,II18845,
    g11659,II18854,g11670,II18857,g11671,II18866,g11682,g11706,g11732,g11734,
    g11735,g11736,g11737,g11740,g11741,g11742,g11743,g11745,g11746,g11747,
    g11748,II18929,g10711,g11749,g11758,g11761,g11762,g11763,g11764,g11765,
    g11766,II18943,g11769,g11770,g11774,g11775,g11776,g11777,g11778,g11779,
    g11782,g11783,II18962,g11786,g11787,II18969,g11791,g11794,g11795,g11796,
    g11797,g11798,g11801,g11802,g11803,g11804,g11808,g11809,II18990,g11812,
    g11813,g11817,g11818,g11819,g11820,g11821,g11824,g11825,g11826,g11827,
    g11829,g11834,g11835,g11836,g11837,g11841,g11842,II19025,g11845,g11846,
    II19030,g11848,g11852,g11853,g11854,g11856,g11857,g11858,g11859,g11862,
    g11866,g11867,g11868,g11869,g11871,g11876,g11877,g11878,g11879,g11883,
    g11884,g11886,g11887,g11888,g11891,g11892,g11893,g11894,g11895,g11898,
    g11899,g11900,g11901,g11904,g11908,g11909,g11910,g11911,g11913,g11918,
    g11919,g11920,g11921,II19105,g11923,g11927,g11929,g11930,g11931,g11932,
    g11933,g11936,II19119,g11937,g11941,g11942,g11943,g11944,g11945,g11948,
    g11949,g11950,g11951,g11954,g11958,g11959,g11960,g11961,g11963,g11968,
    g11969,g11970,g11971,g11972,g11973,II19160,g11976,g11982,g11983,g11984,
    g11985,g11986,g11989,II19174,g11990,g11994,g11995,g11996,g11997,g11998,
    g12001,g12002,g12003,g12004,g12007,II19195,g12009,g12013,g12017,g12020,
    g12021,g12022,g12023,g12024,g12025,II19208,g12027,II19211,g12030,g12037,
    g12038,g12039,g12040,g12041,g12042,II19226,g12045,g12051,g12052,g12053,
    g12054,g12055,g12058,II19240,g12059,g12063,g12064,g12065,g12066,g12067,
    g12071,g12075,g12076,g12077,g12078,g12084,g12085,g12086,g12087,g12088,
    g12089,II19271,g12091,II19274,g12094,g12101,g12102,g12103,g12104,g12105,
    g12106,II19289,g12109,g12115,g12116,g12117,g12118,g12119,g12122,II19303,
    g12123,II19307,g12125,g12130,g12134,g12135,II19315,g12136,II19318,g12139,
    II19321,g12142,g12147,g12148,g12149,g12150,g12156,g12157,g12158,g12159,
    g12160,g12161,II19342,g12163,II19345,g12166,g12173,g12174,g12175,g12176,
    g12177,g12178,II19360,g12181,g12187,g12191,g12196,g12197,II19374,g12198,
    II19377,g12201,II19380,g12204,g12209,g12210,g12211,g12212,g12218,g12219,
    g12220,g12221,g12222,g12223,II19401,g12225,II19404,g12228,g12235,II19412,
    g12239,II19415,g12242,g12246,g12251,g12252,II19426,g12253,II19429,g12256,
    II19432,g12259,g12264,g12265,g12266,g12267,g12275,II19449,g12279,II19452,
    g12282,II19455,g12285,g12289,g12294,g12295,II19466,g12296,II19469,g12299,
    II19472,g12302,g12308,II19479,g12312,II19482,g12315,II19485,g12318,II19488,
    g12321,g12325,g12332,II19500,g12333,II19503,g12336,II19507,g12340,II19510,
    g12343,II19513,g12346,II19516,g12349,g12354,g8381,g12362,II19523,g12363,
    II19526,g12366,II19530,g12370,II19533,g12373,g12378,II19539,g12379,II19542,
    g12382,II19545,g12385,II19549,g12389,II19552,g8430,g12392,g12408,II19557,
    g12409,II19560,g12412,II19563,g12415,g12420,II19569,g12421,g12424,II19573,
    g12425,II19576,g12426,g12430,II19582,g12432,g12434,II19587,g12435,II19591,
    g12437,g12438,II19595,g10810,g12439,II19598,g12440,II19602,g12442,II19605,
    g10797,g12443,II19608,g10831,g12444,II19611,g12445,II19615,g10789,g12447,
    II19618,g10814,g12448,II19621,g10851,g12449,II19624,g12450,II19628,g10784,
    g12452,II19631,g10801,g12453,II19634,g10835,g12454,II19637,g10872,g12455,
    g12456,II19642,g10793,g12460,II19645,g10818,g12461,II19648,g10855,g12462,
    g12463,g12466,II19654,g10805,g12470,II19657,g10839,g12471,g12472,g12473,
    g12476,g12478,g12481,II19667,g10822,g12485,g12490,g12493,g12495,g12498,
    g12502,g12504,g12505,g12510,g12513,g12515,g12518,II19689,g12519,g12521,
    g12522,g12527,g12530,g12532,g12533,II19702,g12534,g12536,g12537,g12542,
    II19711,g12543,g12545,g12546,g12547,II19718,g12548,g12551,II19722,g12552,
    g12553,g12554,II19727,g12555,g12558,g12559,g12560,II19733,g12561,II19736,
    g12564,II19739,g12565,g12596,g12597,g12598,g12599,g12600,II19747,g12601,
    II19750,g12604,II19753,g12607,II19756,g12608,II19759,g12611,g12642,g12643,
    g12644,g12645,g12646,II19767,g12647,II19771,g10038,g12651,II19774,g12654,
    II19777,g12657,g12688,g12689,g12690,g12691,II19784,g12692,II19787,g12695,
    II19791,g12699,II19794,g10676,g12702,II19797,g10147,g12705,II19800,g12708,
    II19803,g12711,g12742,g12743,II19808,g12744,g12748,II19813,g10649,g12749,
    II19816,g10703,g12752,II19820,g12756,II19823,g10705,g12759,II19826,g10252,
    g12762,II19829,g12765,g12768,II19833,g12769,II19836,g12772,g12775,g12776,
    g12782,II19844,g8533,g12783,II19847,g10677,g12786,g12790,II19852,g10679,
    g12791,II19855,g10723,g12794,II19859,g12798,II19862,g10725,g12801,II19865,
    g10354,g12804,g12807,II19869,g12808,II19872,g12811,g12815,II19877,g8547,
    g12816,g12821,II19883,g8550,g12822,II19886,g10706,g12825,g12829,II19891,
    g10708,g12830,II19894,g10744,g12833,II19898,g12837,II19901,g10746,g12840,
    g12843,II19905,g12844,g12847,g12848,g12850,g12851,g12853,II19915,g8560,
    g12854,g12859,II19921,g8563,g12860,II19924,g10726,g12863,g12867,II19929,
    g10728,g12868,II19932,g10763,g12871,g12874,g12875,g12881,g12882,g12891,
    g12892,g12894,II19952,g8571,g12895,g12900,II19958,g8574,g12901,II19961,
    g10747,g12904,g12907,g12909,g12914,g12915,g12921,g12922,g12931,g12932,
    g12934,II19986,g8577,g12935,g12940,g12943,g12944,g12950,g12951,g12960,
    g12961,II20009,g12962,g12965,g12969,g12972,g12973,g12979,g12980,g12993,
    g12996,g12997,g12998,g13003,II20062,g10480,g13011,g13025,g13033,g13036,
    g13043,g13046,g13049,g13057,g13060,g13063,g13066,II20117,g13070,g13073,
    g13076,g13079,g13092,g13095,g13101,g13107,g13117,g13130,g13141,g13148,
    g13151,g13152,g13153,g13154,g13157,g13158,g13159,g13161,g13162,g13163,
    g13166,g13167,g13168,g13169,g13170,g13172,g13173,g13174,g13176,g13177,
    g13178,g13179,g13180,g13181,g13183,g13184,g13185,g13186,g13187,g13188,
    g13189,g13190,g13191,g13192,g13193,g13195,g13196,g13197,g13198,g13199,
    g13200,g13201,g13202,g13203,g13204,g13205,g13206,g13207,g13208,g13209,
    g13210,g13211,g13212,g13213,g13214,II20264,g13215,g13218,g13219,g13220,
    g13221,g13222,g13223,g13224,g13225,g13226,g13227,II20278,g13229,g13232,
    g13233,II20283,g13234,g13237,g13238,g13239,g13240,g13241,g13242,g13243,
    g13244,II20295,g13246,II20299,g13248,g13249,g13250,II20305,g13252,g13255,
    g13256,II20310,g13257,g13260,g13261,g13262,g13263,g13264,g13265,II20320,
    g13267,g13268,II20324,g13269,II20328,g13271,g13272,g13273,II20334,g13275,
    g13278,g13279,II20339,g13280,g13283,g13284,g13285,II20347,g13290,II20351,
    g13292,g13293,II20355,g13294,II20359,g13296,g13297,g13298,II20365,g13300,
    g13303,g13304,g13308,g13309,II20376,g13317,II20379,g13318,II20382,g13319,
    II20386,g13321,II20390,g13323,g13324,II20394,g13325,II20398,g13327,g13328,
    g13329,g13330,II20407,g13336,II20410,g13339,II20414,g13341,II20417,g13342,
    II20421,g13344,II20425,g13346,g13347,g13351,g13352,II20441,g13356,II20444,
    g13359,II20448,g13361,II20451,g13364,II20455,g13366,II20458,g13367,II20462,
    g13369,g13373,II20476,g13381,II20479,g13384,II20483,g13386,II20486,g13389,
    II20490,g13391,II20493,g13394,II20497,g13396,II20500,g13397,g13398,g13400,
    II20514,II20517,II20520,II20523,II20526,II20529,II20532,II20535,II20538,
    II20541,II20544,II20547,II20550,II20553,II20556,II20559,II20562,II20565,
    II20568,II20571,II20574,II20577,II20580,II20583,II20586,II20589,II20592,
    II20595,II20598,II20601,II20604,II20607,II20610,II20613,II20616,II20619,
    II20622,II20625,II20628,II20631,II20634,II20637,II20640,II20643,II20646,
    II20649,II20652,II20655,II20658,II20661,II20664,II20667,II20670,II20673,
    II20676,II20679,II20682,II20685,II20688,II20691,II20694,II20697,II20700,
    II20703,II20706,g13469,II20709,g13519,g13228,g13530,g13251,g13541,g13274,
    g13552,g13299,g13565,g12192,g13568,g11627,II20791,g13149,g13571,II20794,
    g13111,g13572,g13573,g12247,g13576,g11650,II20799,g13155,g13579,II20802,
    g13160,g13580,II20805,g13124,g13581,g13582,g12290,g13585,g11669,II20810,
    g13164,g13588,II20813,g13589,II20816,g12487,g13598,II20820,g13171,g13600,
    II20823,g13135,g13601,g13602,g12326,g13605,g11681,II20828,g13175,g13608,
    II20832,g12507,g13610,II20836,g13182,g13612,II20839,g13143,g13613,g13614,
    g11690,II20844,g12524,g13620,II20848,g13194,g13622,II20852,g12457,g13624,
    g13626,g11697,II20858,g12539,g13632,II20863,g12467,g13635,g13637,g11703,
    g13644,II20873,g12482,g13647,g13649,g11711,g13657,g13669,g13670,II20886,
    g12499,g13673,g13677,g13687,g13699,g13700,g13706,g13714,g13724,g13736,
    g13737,II20909,g13055,g13741,g13750,g13756,g13764,g13774,g13786,g13791,
    g13797,g13805,g13817,g13819,g13825,g13836,g13838,g13840,g13848,g11744,
    g13849,g13850,g13852,g13856,g11759,g13857,g11760,g13858,g13859,g13861,
    II20959,g11713,g13863,g13864,g11767,g13866,g11772,g13867,g11773,g13868,
    g13869,g13872,g11780,g13873,g12698,g13879,g11784,g13881,g11789,g13882,
    g11790,g13883,g13885,g11799,g13886,g12747,g13894,g11806,g13895,g12755,
    g13901,g11810,g13903,g11815,g13906,g11822,g13907,g12781,g13918,g11830,
    g13922,g11831,g13926,g11832,g13927,g12789,g13935,g11839,g13936,g12797,
    g13942,g11843,g13945,g11855,g13946,g12814,II21012,g12503,g13954,g13958,
    g11863,g13962,g11864,g13963,g12820,g13974,g11872,g13978,g11873,g13982,
    g11874,g13983,g12828,g13991,g11881,g13992,g12836,g13999,g11889,g14000,
    g11890,g14001,g12849,II21037,g12486,g14008,g14011,g11896,g14015,g11897,
    g14016,g12852,II21045,g12520,g14024,g14028,g11905,g14032,g11906,g14033,
    g12858,g14044,g11914,g14048,g11915,g14052,g11916,g14053,g12866,g14061,
    g11928,g14062,g12880,II21064,g13147,g14068,g14071,g11934,g14079,g11935,
    g14086,g11938,g14090,g11939,g14091,g11940,g14092,g12890,II21075,g12506,
    g14099,g14102,g11946,g14106,g11947,g14107,g12893,II21083,g12535,g14115,
    g14119,g11955,g14123,g11956,g14124,g12899,g14135,g11964,g14139,g11965,
    II21096,g14144,g14148,g12912,g14153,g12913,g14158,g11974,g14165,g11975,
    g14171,g11979,g14175,g11980,g14176,g11981,g14177,g12920,II21108,g13150,
    g14183,g14186,g11987,g14194,g11988,g14201,g11991,g14205,g11992,g14206,
    g11993,g14207,g12930,II21119,g12523,g14214,g14217,g11999,g14221,g12000,
    g14222,g12933,II21127,g12544,g14230,g14234,g12008,g14238,g12939,g14244,
    g12026,g14249,g12034,g14252,g12035,g14256,g12036,II21137,g14259,g14263,
    g12941,g14268,g12942,g14273,g12043,g14280,g12044,g14286,g12048,g14290,
    g12049,g14291,g12050,g14292,g12949,II21149,g13156,g14298,g14301,g12056,
    g14309,g12057,g14316,g12060,g14320,g12061,g14321,g12062,g14322,g12959,
    II21160,g12538,g14329,g14332,g12068,II21165,g13110,g14337,g14342,g12967,
    g14347,g12079,g14352,g12081,g14355,g12082,g14359,g12083,g14360,g12968,
    g14366,g12090,g14371,g12098,g14374,g12099,g14378,g12100,II21178,g14381,
    g14385,g12970,g14390,g12971,g14395,g12107,g14402,g12108,g14408,g12112,
    g14412,g12113,g14413,g12114,g14414,g12978,II21190,g13165,g14420,g14423,
    g12120,g14431,g12121,g14438,g12124,g14442,g11768,g14450,g12146,g14454,
    g12991,g14459,g12151,g14464,g12153,g14467,g12154,g14471,g12155,g14472,
    g12992,g14478,g12162,g14483,g12170,g14486,g12171,g14490,g12172,II21208,
    g14493,g14497,g12994,g14502,g12995,g14507,g12179,g14514,g12180,g14520,
    g12184,g14524,g12185,g14525,g12195,g14529,g11785,g14537,g12208,g14541,
    g13001,g14546,g12213,g14551,g12215,g14554,g12216,g14558,g12217,g14559,
    g13002,g14565,g12224,g14570,g12232,g14573,g12233,g14577,g12234,g14580,
    g12250,g14584,g11811,g14592,g12263,g14596,g13022,g14601,g12268,g14606,
    g12270,g14609,g12271,g14613,g12272,g14614,g12293,g14618,g11844,g14626,
    g12306,II21241,g13378,g14630,g14637,g12329,g14641,g11823,II21246,g11624,
    g14642,II21249,g11600,g14650,II21252,g11644,g14657,g14668,g11865,II21256,
    g11647,g14669,II21259,g11630,g14677,II21262,g14684,g14685,g12245,II21267,
    g11663,g14691,g14702,g11907,II21271,g11666,g14703,II21274,g11653,g14711,
    II21277,g14718,g14719,g12288,II21282,g11675,g14725,g14736,g11957,II21286,
    g11678,g14737,II21289,g14745,II21292,g14746,g14747,g12324,II21297,g11687,
    g14753,g14764,II21301,g14765,II21304,g14766,g14768,g12352,II21310,g14774,
    II21313,g14775,g14776,g12033,g14794,II21318,g14795,II21321,g14796,g14797,
    g12080,g14811,g12097,II21326,g14829,II21329,g14830,g14831,g11828,g14837,
    g12145,g14849,g12152,g14863,g12169,g14881,II21337,g14882,II21340,g14883,
    g14885,g11860,g14895,g12193,g14904,g11870,g14910,g12207,g14922,g12214,
    g14936,g12231,II21351,g14954,II21354,g14955,g14959,II21361,g13026,g14960,
    II21364,g13028,g14963,g14966,g11902,g14976,g12248,g14985,g11912,g14991,
    g12262,g15003,g12269,g15017,II21374,g15018,II21377,g15019,II21381,g15021,
    g15022,g11781,g15032,g15033,II21389,g12883,g15034,II21392,g13020,g15037,
    II21395,g13034,g15040,II21398,g13021,g15043,g15048,II21404,g13037,g15049,
    II21407,g13039,g15052,g15055,g11952,g15065,g12291,g15074,g11962,g15080,
    g12305,II21415,g15092,II21420,g15095,g15096,g11800,II21426,g11661,g15106,
    II21429,g13027,g15109,II21432,g13044,g15112,II21435,g11662,g15115,g15118,
    g11807,g15128,g15129,II21443,g12923,g15130,II21446,g13029,g15133,II21449,
    g13047,g15136,II21452,g13030,g15139,g15144,II21458,g13050,g15145,II21461,
    g13052,g15148,g15151,g12005,g15161,g12327,g15170,g15174,g15175,g15176,
    g15177,g12339,II21476,g11672,g15179,II21479,g13035,g15182,II21482,g13058,
    g15185,g15188,g11833,II21488,g11673,g15198,II21491,g13038,g15201,II21494,
    g13061,g15204,II21497,g11674,g15207,g15210,g11840,g15220,g15221,II21505,
    g12952,g15222,II21508,g13040,g15225,II21511,g13064,g15228,II21514,g13041,
    g15231,g15236,II21520,g13067,g15237,II21523,g13069,g15240,II21531,g11683,
    g15248,II21534,g13045,g15251,II21537,g13071,g15254,g15260,g15261,g15262,
    g15263,g12369,II21548,g11684,g15265,II21551,g13048,g15268,II21554,g13074,
    g15271,g15274,g11875,II21560,g11685,g15284,II21563,g13051,g15287,II21566,
    g13077,g15290,II21569,g11686,g15293,g15296,g11882,g15306,g15307,II21577,
    g12981,g15308,II21580,g13053,g15311,II21583,g13080,g15314,II21586,g13054,
    g15317,g15322,g15323,II21595,g11691,g15326,II21598,g13059,g15329,II21601,
    g13087,g15332,II21609,g11692,g15340,II21612,g13062,g15343,II21615,g13090,
    g15346,g15352,g15353,g15354,g15355,g12388,II21626,g11693,g15357,II21629,
    g13065,g15360,II21632,g13093,g15363,g15366,g11917,II21638,g11694,g15376,
    II21641,g13068,g15379,II21644,g13096,g15382,II21647,g11695,g15385,g15390,
    II21655,g11696,g15393,II21658,g13072,g15396,II21661,g13098,g15399,II21666,
    g13100,g15404,g15408,g15409,II21674,g11698,g15412,II21677,g13075,g15415,
    II21680,g13102,g15418,II21688,g11699,g15426,II21691,g13078,g15429,II21694,
    g13105,g15432,g15438,g15439,g15440,g15441,g12418,II21705,g11700,g15443,
    II21708,g13081,g15446,II21711,g13108,g15449,g15458,II21720,g11701,g15461,
    II21723,g13088,g15464,II21726,g13112,g15467,II21730,g13089,g15471,g15474,
    II21736,g11702,g15477,II21739,g13091,g15480,II21742,g13114,g15483,II21747,
    g13116,g15488,g15492,g15493,II21755,g11704,g15496,II21758,g13094,g15499,
    II21761,g13118,g15502,II21769,g11705,g15510,II21772,g13097,g15513,II21775,
    g13121,g15516,II21780,g13305,g15521,g15524,g15525,II21787,g11707,g15528,
    II21790,g13099,g15531,II21793,g13123,g15534,II21796,g11708,g15537,g15544,
    II21803,g11709,g15547,II21806,g13103,g15550,II21809,g13125,g15553,II21813,
    g13104,g15557,g15560,II21819,g11710,g15563,II21822,g13106,g15566,II21825,
    g13127,g15569,II21830,g13129,g15574,g15578,g15579,II21838,g11712,g15582,
    II21841,g13109,g15585,II21844,g13131,g15588,II21852,g11716,g15596,II21855,
    g13113,g15599,g15602,g15603,II21862,g11717,g15606,II21865,g13115,g15609,
    II21868,g13134,g15612,II21871,g11718,g15615,g15622,II21878,g11719,g15625,
    II21881,g13119,g15628,II21884,g13136,g15631,II21888,g13120,g15635,g15638,
    II21894,g11720,g15641,II21897,g13122,g15644,II21900,g13138,g15647,II21905,
    g13140,g15652,II21908,g13082,g15655,g15659,g15665,II21918,g11721,g15667,
    II21923,g11722,g15672,II21926,g13126,g15675,g15678,g15679,II21933,g11723,
    g15682,II21936,g13128,g15685,II21939,g13142,g15688,II21942,g11724,g15691,
    g15698,II21949,g11725,g15701,II21952,g13132,g15704,II21955,g13144,g15707,
    II21959,g13133,g15711,II21962,g13004,g15714,g15722,g15724,II21974,g11726,
    g15726,II21979,g11727,g15731,II21982,g13137,g15734,g15737,g15738,II21989,
    g11728,g15741,II21992,g13139,g15744,II21995,g13146,g15747,II21998,g11729,
    g15750,g15762,g15764,II22014,g11730,g15766,II22019,g11731,g15771,II22022,
    g13145,g15774,II22025,g11617,g15777,g15790,g15792,II22044,g11733,g15794,
    g15800,g15813,g15859,II22120,g15876,g15880,g15890,g15904,g15913,g15923,
    g15933,g15942,g15952,g15962,g15971,g15981,II22163,g12433,g15989,g15991,
    g15994,g15997,g16001,g16002,g16005,g16007,g16011,g16012,g16013,g16014,
    g16023,g16024,g16025,g16026,g16027,g16034,g16035,g16039,g16040,g16041,
    g16042,g16043,g16044,g16054,g16055,g16056,g16057,g16061,g16062,g16063,
    g16064,g16065,g16075,g11861,g16088,g16090,g16091,g16092,g16093,g16097,
    g16098,g16099,g16113,g11903,g16126,g16128,g16129,g16130,g16131,g16142,
    g16154,g12194,g16164,g11953,g16177,g16179,g16180,g16189,g16201,g16213,
    g12249,g16223,g12006,g16236,g16243,g16254,g16266,g16278,g12292,g16287,
    g16293,II22382,g16302,g16313,g16325,g16337,g12328,g16351,II22414,g16360,
    g16371,g16395,II22444,g16404,g16433,II22475,g16466,II22503,II22506,II22509,
    II22512,II22515,II22518,II22521,II22524,II22527,II22530,II22533,II22536,
    II22539,II22542,II22545,II22548,II22551,II22554,II22557,II22560,II22563,
    II22566,II22569,II22572,II22575,II22578,II22581,II22584,II22587,II22590,
    II22593,g16501,II22599,g16506,g16507,II22604,g16514,g16515,g16523,II22611,
    g16528,g16529,II22618,g16540,g16543,g16546,g16554,II22626,g16559,g16560,
    II22640,g16572,g16575,g16578,g16586,II22651,g16596,g16599,g16602,II22657,
    g16608,II22663,g16616,g16619,II22667,g16622,II22671,g16626,II22676,g16633,
    II22679,g16636,II22683,g16640,II22687,g16644,II22690,g16647,II22694,g16651,
    II22699,g16656,II22702,g16659,g16665,II22715,g16673,II22718,g16676,g16682,
    g16686,II22726,g16694,g16697,II22730,g16702,g16708,g16712,II22737,g16719,
    g16722,II22741,g16725,g16728,II22745,g16733,g16739,g16743,g16749,g15782,
    II22752,g16758,II22755,g16761,g16764,II22759,g16767,g16770,II22763,g16775,
    g16781,II22768,g16785,II22771,g16788,g16791,II22775,g16794,g16797,g16804,
    g15803,g16809,g15842,II22783,g16813,II22786,g16814,II22789,g16817,g16820,
    g16825,g15855,II22797,g16830,II22800,g16831,II22803,g16832,g16836,g15818,
    g16840,g15878,II22810,g16842,II22813,g16843,g16846,g15903,II22820,g16848,
    II22823,g16849,II22828,g16852,II22836,g16858,II22842,g16862,II22845,g16863,
    g16867,II22852,g16877,II22855,g16878,II22860,g16881,g16884,g16895,II22866,
    g16905,II22869,g16906,II22875,g16910,g16913,g16924,II22881,g16934,II22893,
    g16940,g16943,g16954,II22912,g16971,g16974,g17029,g17057,g17063,g17092,
    g17098,g17130,g17136,g17157,II23253,g17189,II23274,g17200,g17203,II23287,
    g17207,g17208,II23292,g17212,g17214,g17217,II23309,g16132,g17227,II23314,
    g15720,g17230,II23317,g16181,g17233,II23323,g15664,g17237,II23326,g15758,
    g17240,II23329,g15760,g17243,II23335,g16412,g17249,II23338,g15721,g17252,
    II23341,g15784,g17255,g17258,g16053,II23345,g15723,g17259,II23348,g15786,
    g17262,II23351,g15788,g17265,II23358,g16442,g17272,II23361,g15759,g17275,
    II23364,g15805,g17278,g17281,g16081,II23368,g16446,g17282,II23371,g15761,
    g17285,II23374,g15807,g17288,II23377,g15763,g17291,II23380,g15809,g17294,
    II23383,g15811,g17297,II23386,g17300,II23392,g13476,g17304,II23395,g15785,
    g17307,II23398,g15820,g17310,g17313,g16109,g17314,g16110,II23403,g13478,
    g17315,II23406,g15787,g17318,II23409,g15822,g17321,II23412,g13482,g17324,
    II23415,g15789,g17327,II23418,g15824,g17330,II23421,g15791,g17333,II23424,
    g15826,g17336,II23430,g13494,g17342,II23433,g15806,g17345,II23436,g15832,
    g17348,g17351,g16152,II23442,g13495,g17354,II23445,g15808,g17357,II23448,
    g15834,g17360,II23451,g13497,g17363,II23454,g15810,g17366,II23457,g15836,
    g17369,II23460,g13501,g17372,II23463,g15812,g17375,II23466,g15838,g17378,
    II23472,g13510,g17384,II23475,g15821,g17387,II23478,g15844,g17390,g17394,
    g16197,II23487,g13511,g17399,II23490,g15823,g17402,II23493,g15846,g17405,
    II23498,g13512,g17410,II23501,g15825,g17413,II23504,g15848,g17416,II23507,
    g13514,g17419,II23510,g15827,g17422,II23513,g15850,g17425,II23518,g15856,
    g17430,II23521,g13518,g17433,II23524,g15833,g17436,II23527,g15858,g17439,
    II23530,g17442,g17445,g16250,II23539,g13524,g17451,II23542,g15835,g17454,
    II23545,g15867,g17457,II23553,g13525,g17465,II23556,g15837,g17468,II23559,
    g15869,g17471,II23564,g13526,g17476,II23567,g15839,g17479,II23570,g15871,
    g17482,II23575,g15843,g17487,II23578,g15879,g17490,II23581,g13528,g17493,
    II23584,g15845,g17496,g17499,g16292,II23588,g17500,II23591,g17503,II23599,
    g15887,g17511,II23602,g13529,g17514,II23605,g15847,g17517,II23608,g15889,
    g17520,II23611,g17523,II23619,g13535,g17531,II23622,g15849,g17534,II23625,
    g15898,g17537,II23633,g13536,g17545,II23636,g15851,g17548,II23639,g15900,
    g17551,II23645,g13537,g17557,II23648,g15857,g17560,II23651,g13538,g17563,
    g17566,g16346,II23655,g17567,II23658,g17570,II23661,g16085,g17573,II23667,
    g15866,g17579,II23670,g15912,g17582,II23673,g13539,g17585,II23676,g15868,
    g17588,II23679,g17591,II23682,g17594,II23689,g15920,g17601,II23692,g13540,
    g17604,II23695,g15870,g17607,II23698,g15922,g17610,II23701,g17613,II23709,
    g13546,g17621,II23712,g15872,g17624,II23715,g15931,g17627,II23725,g13547,
    g17637,g17640,II23729,g17645,g17648,g16384,II23733,g17649,II23739,g13548,
    g17655,II23742,g15888,g17658,II23745,g13549,g17661,II23748,g17664,II23751,
    g17667,II23754,g16123,g17670,II23760,g15897,g17676,II23763,g15941,g17679,
    II23766,g13550,g17682,II23769,g15899,g17685,II23772,g17688,II23775,g17691,
    II23782,g15949,g17698,II23785,g13551,g17701,II23788,g15901,g17704,II23791,
    g15951,g17707,II23794,g17710,g17720,g15853,g17724,II23817,g13557,g17738,
    g17741,II23821,g17746,II23824,g17749,II23830,g13558,g17755,II23833,g15921,
    g17758,II23836,g13559,g17761,II23839,g17764,II23842,g17767,II23845,g16174,
    g17770,II23851,g15930,g17776,II23854,g15970,g17779,II23857,g13560,g17782,
    II23860,g15932,g17785,II23863,g17788,II23866,g17791,II23874,g15797,g17799,
    g17802,II23888,g17815,g17825,II23904,g13561,g17839,g17842,II23908,g17847,
    II23911,g17850,II23917,g13562,g17856,II23920,g15950,g17859,II23923,g13563,
    g17862,II23926,g17865,II23929,g17868,II23932,g16233,g17871,g17878,g15830,
    g17882,g17892,g17893,II23954,g17903,g17914,II23976,g17927,g17937,II23992,
    g13564,g17951,g17954,II23996,g17959,II23999,g17962,g17969,g15841,g17974,
    g17984,g17988,g17991,g17993,g18003,g18004,II24049,g18014,g18025,II24071,
    g18038,g18048,g18063,g15660,g18070,g15854,g18074,g18084,g18089,g18091,
    g18101,g18105,g18108,g18110,g18120,g18121,II24144,g18131,g18142,II24166,
    g18155,II24171,g16439,g18166,g18170,g15877,g18174,g18179,g18188,g18190,
    g18200,g18205,g18207,g18217,g18221,g18224,g18226,g18236,g18237,II24247,
    g18247,II24258,g16463,g18258,g18261,g15719,g18265,g18275,II24285,g15992,
    g18278,g18281,g18286,g18295,g18297,g18307,g18312,g18314,g18324,g18328,
    g18331,II24346,g15873,g18334,g18337,g15757,g18341,g18351,g18353,II24368,
    g15990,g18355,g18358,g18368,II24394,g15995,g18371,g18374,g18379,g18388,
    g18390,g18400,g18405,g18407,g15959,g18414,g15718,g18415,g15783,g18429,
    II24459,g13599,g18432,g18435,g18436,g18446,g18448,II24481,g15993,g18450,
    g18453,g18463,II24507,g15999,g18466,g18469,g18474,g18483,g18485,g15756,
    g18486,g15804,g18490,g18502,II24560,g13611,g18505,g18508,g18509,g18519,
    g18521,II24582,g15996,g18523,g18526,g18536,II24608,g16006,g18539,g18543,
    g15819,g18552,g18554,g18566,II24662,g13621,g18569,g18572,g18573,g18583,
    g18585,II24684,g16000,g18587,g18593,g15831,g18602,g18604,g18616,II24732,
    g13633,g18619,g18622,g18634,g18636,g18643,g18646,g16341,g18656,g18670,
    g18679,g18691,g18692,g18699,g18708,g18720,g18725,g13865,g18727,g18728,
    g18735,g18744,g18756,g18757,g18758,g18764,g18765,g18772,g18783,g18784,
    g18785,g18786,g18787,g18788,g18789,g18795,g18796,g18805,g18806,g18807,
    g18808,g18809,g18810,g18811,g18812,g18813,g18814,g18815,g18822,g18823,
    g18824,g18825,g18826,g18827,g18828,g18829,g18830,g18831,g18832,g18833,
    g18834,g18838,g18839,g18840,g18841,g18842,g18843,g18844,g18845,g18846,
    g18847,g18848,g18849,g18850,g18851,g18853,g18854,g18855,g18856,g18857,
    g18858,g18859,g18860,g18861,g18862,g18863,g18864,g18865,II24894,g18869,
    g18870,g18871,g18872,g18873,g18874,g18875,g18876,g18877,g18878,g18879,
    g18880,g18881,g18882,g18884,II24913,g18886,II24916,g18890,g18891,g18892,
    g18893,g18894,II24923,g18895,g18896,g18897,g18898,g18899,g18900,g18901,
    g18902,g18903,g18904,g18905,g18908,g18909,g18910,g18911,g18912,II24943,
    g18913,g18914,g18915,g18916,g18917,II24950,g18918,g18919,g18920,g18921,
    g18922,g18923,g18924,g18925,g18926,g18927,g18928,g18929,g18930,g18931,
    II24966,g18932,g18933,g18934,g18935,g18936,II24973,g18937,g18938,g18939,
    g18940,g18941,g18943,II24982,g18944,g18945,g18946,g18947,g18948,g18949,
    g18950,g18951,II24992,g18952,g18953,g18954,g18955,g18956,g18958,II25001,
    g18959,II25004,g18960,g18961,g18962,g18963,g18964,g18965,g18966,g18967,
    II25015,g18969,II25018,g18970,II25021,g18971,g18972,g18973,g18974,g18976,
    II25037,g18981,II25041,g18983,II25044,g18984,II25047,g18985,II25050,g18986,
    g18987,II25054,g18988,II25057,g18989,II25061,g18991,II25064,g18992,II25067,
    g18993,II25071,g18995,II25074,g18996,II25078,g18998,II25081,g18999,II25084,
    g19000,g19001,II25089,g19008,II25092,g19009,II25096,g19011,II25099,II25102,
    II25105,II25108,II25111,II25114,II25117,II25120,II25123,II25126,II25129,
    II25132,II25135,II25138,II25141,II25144,II25147,II25150,II25153,II25156,
    II25159,II25162,II25165,II25168,II25171,II25174,II25177,II25180,II25183,
    II25186,II25189,II25192,II25195,II25198,II25201,II25204,II25207,II25210,
    II25213,II25216,II25219,II25222,II25225,II25228,II25231,II25234,II25237,
    II25240,II25243,II25246,II25249,II25253,g17124,g19064,g19070,II25258,
    g19075,g19078,II25264,g17151,g19081,II25272,g17051,g19091,g19096,g18980,
    II25283,g17086,g19098,II25294,g19105,II25303,g19110,II25308,g19113,II25315,
    g19118,II25320,g19125,II25325,g19132,II25334,g19145,II25338,g19147,II25344,
    g19151,II25351,g19156,II25355,g18669,g19158,II25358,g18678,g19159,II25365,
    g18707,g19164,II25371,g18719,g19168,II25374,g18726,g19169,II25377,g18743,
    g19170,II25383,g18755,g19174,II25386,g18763,g19175,II25389,g18780,g19176,
    II25395,g18782,g19180,II25399,g18794,g19182,II25402,g18821,g19183,II25406,
    g18804,g19185,II25412,g18820,g19189,II25415,g18835,g19190,II25423,g18852,
    g19196,II25426,g18836,g19197,II25429,g18975,g19198,II25432,g18837,g19199,
    II25442,g18866,g19207,II25445,g18968,g19208,II25456,g18883,g19217,II25459,
    g18867,g19218,II25463,g18868,g19220,II25474,g18885,g19229,II25486,g18754,
    g19237,II25489,g18906,g19238,II25492,g18907,g19239,II25506,g18781,g19247,
    II25510,g18542,g19249,g19251,II25525,g18803,g19258,II25528,g18942,g19259,
    g19265,II25557,g18957,g19270,II25567,g17186,g19272,g19280,g19287,II25612,
    g17197,g19291,g19299,g19301,g19302,g17025,g19305,II25660,g17204,g19309,
    g19319,g19322,g19323,g17059,g19326,II25717,g17209,g19330,II25728,g17118,
    g19335,g19346,g19349,g19350,g17094,g19353,II25768,g17139,g19358,II25778,
    g17145,g19369,g19380,g19383,g19384,g17132,g19387,g16567,g19388,II25816,
    g17162,g19390,II25826,g17168,g19401,g19412,g19415,g19417,g16591,g19418,
    II25862,g17177,g19420,II25872,g17183,g19431,g19441,g17213,g19444,g17985,
    g19448,g19452,g19454,g16611,g19455,II25904,g17194,g19457,g19467,g19468,
    g17216,g19471,g18102,g19475,g19479,g19481,g16629,g19482,g19483,g19484,
    g19490,g19491,g17219,g19494,g18218,g19498,g19502,g19504,g19505,g19511,
    g19512,g17221,g19515,g18325,g19519,g19523,g19524,g19530,g19533,g19534,
    II25966,g16654,g19543,II25971,g16671,g19546,II25977,g16692,g19550,II25985,
    g16718,g19556,II25994,g16860,g19563,II26006,g16866,g19573,g19577,g19578,
    II26025,g16803,g19595,II26028,g16566,g19596,g19607,g19608,II26051,g16824,
    g19622,g19640,g19641,II26078,g16835,g19652,II26085,g18085,g19657,g19680,
    g19681,II26112,g16844,g19689,II26115,g16845,g19690,II26123,g19696,II26134,
    g18201,g19705,II26154,g16851,g19725,II26171,g19740,II26182,g18308,g19749,
    II26195,g16853,g19762,II26198,g16854,g19763,II26220,g19783,II26231,g18401,
    g19792,II26237,g16857,g19798,II26266,g19825,g19830,II26276,g16861,g19838,
    II26334,g18977,g19890,II26337,g16880,g19893,II26340,g19894,II26365,g18626,
    g19915,g19918,II26369,g19919,g19933,g18548,II26388,g19934,II26401,g17012,
    g19945,g19948,g17896,g19950,g18598,II26407,g19951,II26413,g16643,g19957,
    II26420,g17042,g19972,g19975,g18007,g19977,g18630,II26426,g16536,g19978,
    II26437,g16655,g19987,II26444,g17076,g20002,g20005,g18124,g20007,g18639,
    II26458,g20016,II26469,g16672,g20025,II26476,g17111,g20040,g20043,g18240,
    II26481,g18590,g20045,II26494,g20058,II26505,g16693,g20067,II26512,g16802,
    g20082,g20083,g17968,II26535,g20099,II26545,g16823,g20105,II26574,g20124,
    g20127,g18623,g20140,g20163,g17973,II26612,g20164,g20178,g20193,II26642,
    g20198,g20212,g20223,II26664,g20228,g20242,g20250,II26679,g20255,g20269,
    g20273,g20278,g20279,g20281,g20286,g20287,g20288,g20289,g20290,g20292,
    II26714,g20295,g20296,g20297,g20298,g20302,g20303,g20304,g20305,g20306,
    g20308,g20311,g20312,g20313,g20315,g20316,g20317,g20321,g20322,g20323,
    g20324,g20325,g20327,g20328,g20329,g20330,g20331,g20332,g20334,g20335,
    g20336,g20340,g20341,g20342,g20344,g20345,g20346,g20347,g20348,g20349,
    g20350,g20351,g20352,g20354,g20355,g20356,II26777,g17222,g20360,g20361,
    g20362,g20363,g20364,g20365,g20366,g20367,g20368,g20369,g20370,g20371,
    g20372,g20373,g20374,II26796,g17224,g20377,g20378,g20379,g20380,g20381,
    g20382,g20383,g20384,g20385,g20386,g20387,g20388,g20389,g20390,g20391,
    g20392,g20393,g20394,II26816,g17225,g20395,II26819,g17226,g20396,g20397,
    g20398,g20399,g20400,g20401,g20402,g20403,g20404,g20405,g20406,g20407,
    g20408,g20409,g20410,g20411,g20412,g20413,g20414,g20415,g20416,II26843,
    g17228,g20418,II26846,g17229,g20419,g20420,g20421,g20422,g20423,g20424,
    g20425,g20426,g20427,g20428,g20429,g20430,g20431,g20432,g20433,g20434,
    g20435,g20436,g20437,g20438,II26868,g17234,g20439,II26871,g17235,g20440,
    II26874,g17236,g20441,g20442,g20443,g20444,g20445,g20446,g20447,g20448,
    g20449,g20450,g20451,g20452,g20453,g20454,g20455,g20456,II26892,g17246,
    g20457,II26895,g17247,g20458,II26898,g17248,g20459,g20461,g20462,g20463,
    g20464,g20465,g20466,g20467,g20468,II26910,g17269,g20469,II26913,g17270,
    g20470,II26916,g17271,g20471,g20476,g20477,II26923,g17302,g20478,II26926,
    g17303,g20479,II26931,g17340,g20484,II26934,g17341,g20485,g20490,II26940,
    g17383,g20491,g20496,II26947,g17429,g20498,g20500,g20501,g20504,g20505,
    g20507,II26960,g20513,g20516,g20517,g20518,II26966,g20519,g20526,II26972,
    g20531,g20534,g20535,g20536,II26980,g20539,g20545,II26985,g20550,g20553,
    g20554,II26990,II26993,II26996,II26999,II27002,II27005,II27008,II27011,
    II27014,II27017,II27020,II27023,II27026,II27029,II27032,II27035,II27038,
    II27041,II27044,II27047,II27050,II27053,II27056,II27059,II27062,II27065,
    II27068,II27071,II27074,II27077,II27080,II27083,II27086,II27089,II27092,
    II27095,II27098,II27101,II27104,II27107,II27110,II27113,II27116,II27119,
    II27122,II27125,II27128,II27131,II27134,II27137,II27140,II27143,II27146,
    II27149,II27152,II27155,II27158,II27161,II27164,II27167,II27170,II27173,
    II27176,II27179,II27182,II27185,II27188,II27191,II27194,II27197,II27200,
    II27203,II27206,II27209,II27212,II27215,II27218,II27221,II27225,g20634,
    II27228,g20637,II27232,g20641,II27235,g20644,II27240,g20649,II27243,g20652,
    II27246,g20655,II27250,g20659,II27253,g20662,II27257,g20666,II27260,g20669,
    II27264,g20673,II27267,g20676,II27270,g20679,II27275,g20684,II27278,g20687,
    II27281,g20690,II27285,g20694,II27288,g20697,II27293,g20704,II27297,g20708,
    II27300,g20711,II27303,g20714,II27308,g20719,II27311,g20722,II27314,g20725,
    II27318,g20729,II27321,g20732,II27324,g20735,II27328,g20739,II27332,g20743,
    II27335,g20746,II27338,g20749,II27343,g20754,II27346,g20757,II27349,g20760,
    II27352,g20763,II27355,g20766,II27358,g20769,II27361,g20772,II27365,g20776,
    II27369,g20780,II27372,g20783,II27375,g20786,II27379,g20790,II27382,g20793,
    II27385,g20796,II27388,g20799,II27391,g20802,II27395,g20806,II27399,g20810,
    II27402,g20813,II27405,g20816,II27408,g20819,II27411,g20822,II27416,g20827,
    II27419,g20830,II27422,g20833,II27426,g20837,g20842,g20850,g20858,g20866,
    g20885,g19865,g20904,g19896,g20928,g19921,II27488,g20310,g20942,II27491,
    g20314,g20943,g20956,g19936,II27516,g20333,g20971,II27531,g20343,g20984,
    II27534,g20985,II27537,g20986,II27549,g20353,g20998,II27565,g21012,II27577,
    g20375,g21024,II27585,g20376,g21030,II27593,g21036,g21050,II27614,g21057,
    II27621,g20417,g21064,g21066,g21069,g21076,g21079,II27646,g21087,g21090,
    g21093,II27658,g21099,g21102,II27667,g21108,II27672,g21113,II27684,g21125,
    II27689,g21130,II27705,g21144,II27727,g21164,II27749,g19954,g21184,g21187,
    II27766,g19984,g21199,g21202,II27779,g20022,g21214,g21217,II27785,g20064,
    g21222,g21225,g21241,g21249,g21258,g21266,II27822,g21271,II27827,g21278,
    II27832,g21285,II27838,g21293,II27868,g19144,g21327,II27897,g19149,g21358,
    II27900,g21359,II27917,g19153,g21376,II27920,g19154,g21377,II27927,g21382,
    II27942,g19157,g21399,g21400,II27949,g21404,II27958,g21415,II27969,g19162,
    g21426,II27972,g19163,g21427,II27976,g21429,II27984,g21441,II27992,g21449,
    II28000,g19167,g21457,II28003,g21458,g21461,II28009,g20473,g21473,II28013,
    g21477,II28019,g21483,II28027,g21491,II28031,g19172,g21495,II28034,g19173,
    g21496,II28038,g21498,II28043,g21505,g21508,II28047,g20481,g21514,II28051,
    g21518,II28057,g21524,II28061,g19178,g21528,g21529,II28065,g21530,II28072,
    g21537,II28076,g21541,g21544,II28080,g20487,g21550,II28084,g21554,II28087,
    g19184,g21557,II28090,g20008,g21558,II28093,g21561,g21565,II28100,g21566,
    II28107,g21573,II28111,g21577,g21580,II28115,g20493,g21586,II28119,g21590,
    II28123,g21594,g21598,II28130,g21599,II28137,g21606,II28143,g21612,II28148,
    g21619,II28152,g21623,g21627,II28159,g21628,II28169,g21640,II28174,g21647,
    II28178,g21651,II28184,g19103,g21655,g21661,II28201,g21671,II28206,g21678,
    II28210,g20537,g21682,g21690,II28229,g21700,II28235,g20153,g21708,g21716,
    g21726,g21742,g21752,g21766,g21782,II28314,g19152,g21795,II28357,g20497,
    g21824,II28360,g21825,g21861,g21867,g21872,g21876,g21883,g21886,g21895,
    g21902,g21907,II28432,g21914,II28435,g21917,g21921,g21927,II28443,g21928,
    II28447,g21932,II28450,g21935,g21939,II28455,II28458,II28461,II28464,
    II28467,II28470,II28473,II28476,II28479,II28482,II28485,II28488,II28491,
    II28494,II28497,II28500,II28503,II28506,II28509,II28512,II28515,II28518,
    II28521,II28524,II28527,g21407,g21967,II28541,g21467,g21982,II28550,g21432,
    g21995,II28557,g22003,II28564,g21385,g22014,II28628,g21842,g22082,II28649,
    g21843,g22107,II28671,g21845,g22133,II28693,g21847,g22156,II28712,g21851,
    g22176,g22212,g22213,g22217,II28781,g21331,g22219,g22221,g22222,II28789,
    g21878,g22225,II28792,g21880,g22226,g22230,II28800,g21316,g22232,g22233,
    g22236,g22237,g22239,g22240,g22241,II28813,g21502,g22243,g22246,g22248,
    g22251,g22252,II28825,g21882,g22253,g22256,g22257,g22258,II28833,g21470,
    g22259,g22260,g22261,g22262,g22266,g22268,g22271,g22274,g22275,g22276,
    g22277,g22278,g22279,g22283,g22286,g22287,g22290,g22293,g22294,g22295,
    g22296,g22297,g22298,II28876,g21238,g22300,g22303,g22304,g22306,g22307,
    g22310,g22313,g22314,g22315,g22316,g21149,g22318,g22319,g21228,II28896,
    g21246,g22328,g22331,g22332,g22334,g22335,g22338,g22341,g21169,g22343,
    g22344,g21233,II28913,g21255,g22353,g22356,g22357,g22359,g22360,g22364,
    g21189,g22366,g22367,g21242,II28928,g21263,g22376,g22379,g22380,g22384,
    g21204,g22386,g22387,g21250,g22401,g21533,g22402,g21569,g22403,g21602,
    g22404,g21631,II28949,g21685,g22405,g22408,II28953,g21659,g22409,II28956,
    g21714,g22412,II28959,g21636,g22415,II28962,g21721,g22418,g22421,II28966,
    g20633,g22422,II28969,g21686,g22425,II28972,g21736,g22428,II28975,g21688,
    g22431,II28978,g21740,g22434,II28981,g21667,g22437,II28984,g21747,g22440,
    g22443,II28988,g20874,g22444,II28991,g20648,g22445,II28994,g21715,g22448,
    II28997,g21759,g22451,II29001,g20658,g22455,II29004,g21722,g22458,II29007,
    g21760,g22461,II29010,g21724,g22464,II29013,g21764,g22467,II29016,g21696,
    g22470,II29019,g21771,g22473,g22476,II29023,g20672,g22477,II29026,g21737,
    g22480,II29030,g20683,g22484,II29033,g21741,g22487,II29036,g21775,g22490,
    II29040,g20693,g22494,II29043,g21748,g22497,II29046,g21776,g22500,II29049,
    g21750,g22503,II29052,g21780,g22506,II29055,g21732,g22509,II29058,g20703,
    g22512,II29064,g20875,g22518,II29067,g20876,g22519,II29070,g20707,g22520,
    II29073,g21761,g22523,II29077,g20718,g22527,II29080,g21765,g22530,II29083,
    g21790,g22533,II29087,g20728,g22537,II29090,g21772,g22540,II29093,g21791,
    g22543,g22547,II29098,g20879,g22548,II29101,g20880,g22549,II29104,g20881,
    g22550,II29107,g21435,g22551,II29110,g20738,g22552,II29116,g20882,g22558,
    II29119,g20883,g22559,II29122,g20742,g22560,II29125,g21777,g22563,II29129,
    g20753,g22567,II29132,g21781,g22570,II29135,g21804,g22573,II29142,g20682,
    g22582,II29145,g20891,g22583,II29148,g20892,g22584,II29151,g20893,g22585,
    II29154,g20894,g22586,g22588,II29159,g20896,g22589,II29162,g20897,g22590,
    II29165,g20898,g22591,II29168,g20775,g22592,II29174,g20899,g22598,II29177,
    g20900,g22599,II29180,g20779,g22600,II29183,g21792,g22603,g22609,II29191,
    g20901,g22611,II29194,g20902,g22612,II29197,g20903,g22613,II29203,g20717,
    g22619,II29206,g20910,g22620,II29209,g20911,g22621,II29212,g20912,g22622,
    II29215,g20913,g22623,g22625,II29220,g20915,g22626,II29223,g20916,g22627,
    II29226,g20917,g22628,II29229,g20805,g22629,II29235,g20918,g22635,II29238,
    g20919,g22636,II29243,g20921,g22639,II29246,g20922,g22640,II29249,g20923,
    g22641,II29252,g20924,g22642,g22645,II29259,g20925,g22647,II29262,g20926,
    g22648,II29265,g20927,g22649,II29271,g20752,g22655,II29274,g20934,g22656,
    II29277,g20935,g22657,II29280,g20936,g22658,II29283,g20937,g22659,g22661,
    II29288,g20939,g22662,II29291,g20940,g22663,II29294,g20941,g22664,II29301,
    g20944,g22669,II29304,g20945,g22670,II29307,g20946,g22671,II29310,g20947,
    g22672,II29313,g20948,g22673,II29317,g20949,g22675,II29320,g20950,g22676,
    II29323,g20951,g22677,II29326,g20952,g22678,g22681,II29333,g20953,g22683,
    II29336,g20954,g22684,II29339,g20955,g22685,II29345,g20789,g22691,II29348,
    g20962,g22692,II29351,g20963,g22693,II29354,g20964,g22694,II29357,g20965,
    g22695,II29360,g21796,g22696,II29366,g20966,g22702,II29369,g20967,g22703,
    II29372,g20968,g22704,II29375,g20969,g22705,II29378,g20970,g22706,II29383,
    g20972,g22709,II29386,g20973,g22710,II29389,g20974,g22711,II29392,g20975,
    g22712,II29395,g20976,g22713,II29399,g20977,g22715,II29402,g20978,g22716,
    II29405,g20979,g22717,II29408,g20980,g22718,g22721,II29415,g20981,g22723,
    II29418,g20982,g22724,II29421,g20983,g22725,II29426,g20989,g22728,II29429,
    g20990,g22729,II29432,g20991,g22730,II29435,g20992,g22731,II29439,g20993,
    g22733,II29442,g20994,g22734,II29445,g20995,g22735,II29448,g20996,g22736,
    II29451,g20997,g22737,II29456,g20999,g22740,II29459,g21000,g22741,II29462,
    g21001,g22742,II29465,g21002,g22743,II29468,g21003,g22744,II29472,g21004,
    g22746,II29475,g21005,g22747,II29478,g21006,g22748,II29481,g21007,g22749,
    II29484,g21903,g22750,g22753,II29490,g21009,g22756,II29493,g21010,g22757,
    II29496,g21011,g22758,II29500,g21015,g22760,II29503,g21016,g22761,II29506,
    g21017,g22762,II29509,g21018,g22763,II29513,g21019,g22765,II29516,g21020,
    g22766,II29519,g21021,g22767,II29522,g21022,g22768,II29525,g21023,g22769,
    II29530,g21025,g22772,II29533,g21026,g22773,II29536,g21027,g22774,II29539,
    g21028,g22775,II29542,g21029,g22776,g22777,II29547,g21031,g22785,II29550,
    g21032,g22786,g22787,II29556,g21033,g22790,II29559,g21034,g22791,II29562,
    g21035,g22792,II29566,g21039,g22794,II29569,g21040,g22795,II29572,g21041,
    g22796,II29575,g21042,g22797,II29579,g21043,g22799,II29582,g21044,g22800,
    II29585,g21045,g22801,II29588,g21046,g22802,II29591,g21047,g22803,g22805,
    g21894,g22806,g21615,II29600,g21720,g22812,II29603,g21051,g22824,II29606,
    g21364,g22825,II29610,g21052,g22827,II29613,g21053,g22828,g22829,II29619,
    g21054,g22832,II29622,g21055,g22833,II29625,g21056,g22834,II29629,g21060,
    g22836,II29632,g21061,g22837,II29635,g21062,g22838,II29638,g21063,g22839,
    II29641,g20825,g22840,g22843,g21889,g22847,g21643,II29653,g21746,g22852,
    II29656,g21070,g22864,II29660,g21071,g22866,II29663,g21072,g22867,g22868,
    II29669,g21073,g22871,II29672,g21074,g22872,II29675,g21075,g22873,g22875,
    g21884,g22882,g21674,II29687,g21770,g22887,II29690,g21080,g22899,II29694,
    g21081,g22901,II29697,g21082,g22902,II29700,g20700,g22903,g22907,g21711,
    g22917,g21703,II29712,g21786,g22922,II29715,g21094,g22934,II29724,g22945,
    II29727,g20877,g22948,g22949,g21665,g22954,g21739,g22958,g21694,g22962,
    g21763,g22966,g21730,II29736,g20884,g22970,g22971,g21779,g22975,g21756,
    II29741,g21346,g22979,g22980,g21794,g22986,g22988,g22989,g22991,g22995,
    g22996,g22998,g23001,g23002,g23006,g23007,g23008,g23012,g23015,g23016,
    g23020,g23021,g23024,g23028,g23031,g23032,g23036,g23037,g23038,g23041,
    g23045,g23048,g23049,II29797,g23050,II29802,g23055,g23056,g23057,g23060,
    g23064,II29812,g23065,II29817,g23068,g23069,g23074,g23075,II29827,g23078,
    g23079,g23082,g23087,g23088,II29841,g23094,g23095,g23098,g23103,II29852,
    g23105,g23112,g23115,II29863,g23116,II29872,g23125,II29881,g23134,g23140,
    g23141,g23142,g23143,g23144,g23145,g23146,g23147,II29897,II29900,II29903,
    II29906,II29909,II29912,II29915,II29918,II29921,II29924,II29927,II29930,
    II29933,II29936,II29939,II29942,II29945,II29948,II29951,II29954,II29957,
    II29960,II29963,II29966,II29969,II29972,II29975,II29978,II29981,II29984,
    II29987,II29990,II29993,II29996,II29999,II30002,II30005,II30008,II30011,
    II30014,II30017,II30020,II30023,II30026,II30029,II30032,II30035,II30038,
    II30041,II30044,II30047,II30050,II30053,II30056,II30059,II30062,II30065,
    II30068,II30071,II30074,II30077,II30080,II30083,II30086,II30089,II30092,
    II30095,II30098,II30101,II30104,II30107,II30110,II30113,II30116,II30119,
    II30122,II30125,II30128,II30131,II30134,II30137,II30140,II30143,II30146,
    II30149,II30152,II30155,II30158,II30161,II30164,II30167,II30170,II30173,
    II30176,II30179,II30182,II30185,II30188,II30191,II30194,II30197,II30200,
    II30203,II30206,II30209,II30212,II30215,II30218,II30221,II30224,II30227,
    II30230,II30233,II30236,II30239,II30242,II30245,II30248,II30251,II30254,
    II30257,II30260,II30263,II30266,II30269,II30272,II30275,II30278,II30281,
    II30284,II30287,II30290,II30293,II30296,II30299,II30302,II30305,II30308,
    II30311,II30314,II30317,II30320,II30323,II30326,II30329,II30332,II30335,
    II30338,II30341,II30344,II30347,II30350,II30353,II30356,II30359,II30362,
    II30365,II30368,II30371,II30374,II30377,II30380,II30383,II30386,II30389,
    II30392,II30395,II30398,II30401,II30404,II30407,g23403,g23052,g23410,
    g23071,g23415,g23084,g23420,g23089,g23424,g23100,g23429,g23107,g23435,
    g23120,II30467,g23000,g23438,II30470,g23117,g23439,g23441,g23129,g23444,
    II30476,g22876,g23448,II30480,g23014,g23452,II30483,g23126,g23453,II30486,
    g23022,g23454,II30489,g22911,g23455,II30493,g23030,g23459,II30496,g23137,
    g23460,II30501,g23039,g23463,II30504,g22936,g23464,II30508,g23047,g23468,
    II30511,g21970,g23469,g23470,g22188,II30516,g23058,g23472,II30519,g22942,
    g23473,II30525,g23067,g23481,g23482,g22197,II30531,g23076,g23485,II30536,
    g23081,g23492,g23493,g22203,II30544,g23092,g23500,II30547,g23093,g23501,
    II30552,g23097,g23508,g23509,g22209,II30560,g23110,g23516,II30563,g23111,
    g23517,II30568,g23114,g23524,II30575,g23123,g23531,II30578,g23124,g23532,
    II30586,g23132,g23542,II30589,g23133,g23543,II30594,g22025,g23546,II30598,
    g22027,g23548,II30601,g22028,g23549,II30607,g22029,g23553,II30611,g22030,
    g23555,II30614,g22031,g23556,II30617,g22032,g23557,II30623,g22033,g23561,
    II30626,g22034,g23562,II30632,g22035,g23566,II30636,g22037,g23568,II30639,
    g22038,g23569,II30642,g22039,g23570,II30648,g22040,g23574,II30651,g22041,
    g23575,II30654,g22042,g23576,II30660,g22043,g23580,II30663,g22044,g23581,
    II30669,g22045,g23585,II30673,g22047,g23587,II30676,g22048,g23588,II30679,
    g22049,g23589,II30686,g23136,g23594,II30689,g22054,g23595,II30692,g22055,
    g23596,II30695,g22056,g23597,II30701,g22057,g23601,II30704,g22058,g23602,
    II30707,g22059,g23603,II30713,g22060,g23607,II30716,g22061,g23608,II30722,
    g22063,g23612,II30725,g22064,g23613,II30728,g22065,g23614,II30735,g22066,
    g23619,II30738,g22067,g23620,II30741,g22068,g23621,II30748,g21969,g23626,
    II30751,g22073,g23627,II30754,g22074,g23628,II30757,g22075,g23629,II30763,
    g22076,g23633,II30766,g22077,g23634,II30769,g22078,g23635,II30776,g22079,
    g23640,II30779,g22080,g23641,II30782,g22081,g23642,II30786,g22454,g23644,
    II30797,g22087,g23661,II30800,g22088,g23662,II30803,g22089,g23663,II30810,
    g22090,g23668,II30813,g22091,g23669,II30816,g22092,g23670,II30823,g21972,
    g23675,II30826,g22097,g23676,II30829,g22098,g23677,II30832,g22099,g23678,
    II30838,g22100,g23682,II30841,g22101,g23683,II30844,g22102,g23684,II30847,
    g22103,g23685,II30854,g22104,g23690,II30857,g22105,g23691,II30860,g22106,
    g23692,II30864,g22493,g23694,II30875,g22112,g23711,II30878,g22113,g23712,
    II30881,g22114,g23713,II30888,g22115,g23718,II30891,g22116,g23719,II30894,
    g22117,g23720,II30901,g21974,g23725,II30905,g22122,g23727,II30908,g22123,
    g23728,II30911,g22124,g23729,II30914,g22125,g23730,II30917,g23731,II30922,
    g22126,g23736,II30925,g22127,g23737,II30928,g22128,g23738,II30931,g22129,
    g23739,II30938,g22130,g23744,II30941,g22131,g23745,II30944,g22132,g23746,
    II30948,g22536,g23748,II30959,g22138,g23765,II30962,g22139,g23766,II30965,
    g22140,g23767,II30973,g22141,g23773,II30976,g22142,g23774,II30979,g22143,
    g23775,II30985,g22992,g23779,II30988,g22145,g23782,II30991,g22146,g23783,
    II30994,g22147,g23784,II30997,g22148,g23785,II31000,g23786,II31005,g22149,
    g23791,II31008,g22150,g23792,II31011,g22151,g23793,II31014,g22152,g23794,
    II31021,g22153,g23799,II31024,g22154,g23800,II31027,g22155,g23801,II31031,
    g22576,g23803,II31043,g22161,g23821,II31050,g22162,g23826,II31053,g22163,
    g23827,II31056,g22164,g23828,II31062,g23003,g23832,II31065,g22166,g23835,
    II31068,g22167,g23836,II31071,g22168,g23837,II31074,g22169,g23838,II31077,
    g23839,II31082,g22170,g23844,II31085,g22171,g23845,II31088,g22172,g23846,
    II31091,g22173,g23847,g23853,II31102,g22177,g23856,II31109,g22178,g23861,
    II31112,g22179,g23862,II31115,g22180,g23863,II31121,g23017,g23867,II31124,
    g22182,g23870,II31127,g22183,g23871,II31130,g22184,g23872,II31133,g22185,
    g23873,II31136,g23874,II31141,g23879,II31144,g22935,g23882,g23885,g22062,
    g23887,II31152,g22191,g23890,II31159,g22192,g23895,II31162,g22193,g23896,
    II31165,g22194,g23897,II31171,g23033,g23901,g23905,g22046,g23908,II31181,
    g22200,g23911,II31188,g21989,g23916,g23918,g22036,II31195,g22578,g23923,
    g23940,II31205,g22002,g23943,II31213,g22615,g23955,II31226,g22651,g23984,
    II31232,g22026,g24000,II31235,g22218,g24001,II31244,g22687,g24014,II31250,
    g22953,g24030,II31253,g22231,g24033,II31257,g22234,g24035,g24047,g23023,
    II31266,g22242,g24051,II31270,g22247,g24053,II31274,g22249,g24055,g24060,
    g23040,II31282,g22263,g24064,II31286,g22267,g24066,II31290,g22269,g24068,
    g24073,g23059,II31298,g22280,g24077,II31302,g22284,g24079,g24084,g23077,
    II31310,g22299,g24088,g24094,g22339,g24095,g22362,g24096,g24097,g22382,
    g24098,g24099,g24101,g24102,g24103,g22397,g24104,g24105,g24106,g24107,
    g24108,g24110,g24111,g24112,g24113,g24114,g24115,g22381,g24121,g24122,
    g24123,g24124,g24125,g24127,g24128,g24129,g24130,g24131,g24132,g24133,
    g24134,g22396,g24140,g24141,g24142,g24143,g24144,g24146,g24147,g24148,
    g24149,g24150,g24151,g24152,g24153,g22399,g24159,g24160,g24161,g24162,
    g24163,g24164,g24165,g24166,g24167,g24168,g22400,g24175,g24176,g24177,
    g24180,II31387,g22811,g24183,g24210,g24220,II31417,g24233,II31426,g24240,
    II31436,g24248,g24251,II31445,g24255,II31451,II31454,II31457,II31460,
    II31463,II31466,II31469,II31472,II31475,II31478,II31481,II31484,II31487,
    II31490,II31493,II31496,II31499,II31502,II31505,II31508,II31511,II31514,
    II31517,II31520,II31523,II31526,II31529,II31532,II31535,II31538,II31541,
    II31544,II31547,II31550,II31553,II31556,II31559,II31562,II31565,II31568,
    II31571,II31574,II31577,II31580,II31583,II31586,II31589,II31592,II31595,
    II31598,II31601,II31604,II31607,II31610,II31613,II31616,II31619,II31622,
    II31625,II31628,II31631,II31634,II31637,II31640,II31643,II31646,II31649,
    II31652,II31655,II31658,II31661,II31664,II31667,II31670,II31673,II31676,
    II31679,II31682,II31685,II31688,II31691,II31694,II31697,II31700,II31703,
    II31706,II31709,II31712,II31715,II31718,II31721,II31724,II31727,II31730,
    II31733,II31736,II31739,II31742,II31745,II31748,II31751,II31754,II31757,
    II31760,II31763,II31766,II31769,II31772,II31775,II31778,II31781,II31784,
    II31787,II31790,II31793,II31796,II31799,II31802,II31805,II31808,II31811,
    II31814,II31817,II31820,II31823,II31826,II31829,II31832,II31835,II31838,
    II31841,II31844,II31847,II31850,II31853,II31856,II31859,II31862,II31865,
    II31868,II31871,II31874,II31877,II31880,II31883,II31886,II31889,II31892,
    II31895,II31898,II31901,II31904,II31907,II31910,II31913,II31916,II31919,
    II31922,II31925,II31928,II31931,II31934,II31937,II31940,II31943,II31946,
    II31949,g24482,II32042,g23399,g24518,II32057,g23406,g24531,II32067,g24174,
    g24539,II32074,g23413,g24544,II32081,g24178,g24549,II32085,g24179,g24551,
    II32092,g23418,g24556,II32098,g24181,g24560,II32102,g24182,g24562,II32109,
    g24206,g24567,II32112,g24207,g24568,II32116,g24208,g24570,II32120,g24209,
    g24572,II32126,g24212,g24576,II32129,g24213,g24577,II32133,g24214,g24579,
    II32137,g24215,g24581,II32140,g24216,g24582,II32143,g24218,g24583,II32146,
    g24219,g24584,II32150,g24222,g24586,II32153,g24223,g24587,II32156,g24225,
    g24588,II32159,g24226,g24589,II32164,g24228,g24592,II32167,g24230,g24593,
    II32170,g24231,g24594,II32175,g24235,g24597,II32178,g24237,g24598,II32181,
    g24238,g24599,II32184,g23497,g24600,II32189,g24243,g24605,II32193,g23513,
    g24607,II32198,g24250,g24612,II32203,g23528,g24619,II32210,g23539,g24630,
    g24648,g24668,g24687,g24704,II32248,g23919,II32251,g24735,II32281,g23950,
    g24763,II32320,g23979,g24784,II32365,g24009,g24805,g24815,II32388,g23385,
    g24816,II32419,g24043,g24827,g24834,II32439,g23392,g24835,g24850,II32487,
    g23400,g24851,II32506,g23324,g24856,g24864,II32535,g23407,g24865,II32556,
    g23329,g24872,II32583,g23330,g24879,II32604,g23339,g24886,g24893,g23486,
    II32642,g23348,g24903,g24912,g23495,g24916,g23502,g24929,g23511,g24933,
    g23518,g24939,g23660,g24941,g23526,g24945,g23533,II32704,g23357,g24949,
    g24950,g23710,g24952,g23537,II32716,g23358,g24956,II32719,g23359,g24957,
    g24958,g23478,g24962,g23764,g24969,g23489,g24973,g23819,g24982,g23505,
    g24993,g23521,g25087,g25094,g25095,II32829,g24059,g25103,g25104,g25105,
    II32835,g24072,g25109,g25110,g25111,g25115,g25116,II32844,g25118,II32847,
    g24083,g25119,g25120,II32851,g25121,II32854,g24092,g25122,II32857,g25123,
    II32860,g25124,g25126,II32868,II32871,II32874,II32877,II32880,II32883,
    II32886,II32889,II32892,II32895,II32898,II32901,II32904,II32907,II32910,
    II32913,II32916,II32919,II32922,II32925,II32928,II32931,II32934,II32937,
    II32940,II32943,II32946,II32949,II32952,II32955,II32958,II32961,II32964,
    II32967,II32970,II32973,II32976,II32979,II32982,II32985,II32988,II32991,
    II32994,II32997,II33000,II33003,II33006,II33009,II33013,g25179,II33016,
    g25180,g25274,g25283,g25291,II33128,g24975,g25296,g25301,g25305,g24880,
    II33136,g24986,g25306,g25313,g24868,g25314,g24897,II33145,g24997,g25315,
    g25319,g24857,g25322,g24883,g25323,g24920,II33154,g25005,g25324,II33157,
    g25027,g25327,g25329,g24844,g25330,g24873,g25332,g24900,g25333,g24937,
    g25335,g24832,II33168,g25042,g25336,g25338,g24860,g25339,g24887,g25341,
    g24923,g25347,g24817,g25349,g24848,II33182,g25056,g25350,g25352,g24875,
    g25353,g24904,II33188,g24814,g25354,g25355,g24797,g25361,g24837,g25363,
    g24862,II33198,g25067,g25364,g25366,g24889,g25367,g24676,g25368,g24778,
    II33205,g24833,g25369,g25370,g24820,g25376,g24852,g25378,g24877,g25379,
    g25383,g24766,g25384,g24695,g25385,g24801,II33219,g24849,g25386,g25387,
    g24839,g25393,g24866,g25394,g24753,g25395,g25399,g24787,g25400,g24712,
    g25401,g24823,II33232,g24863,g25402,g25403,g24854,g25404,g24771,g25405,
    g25409,g24808,g25410,g24723,g25411,g24842,g25412,g24791,g25413,g25417,
    g24830,g25419,g24812,II33246,g24890,II33249,g25421,g25422,g25430,g24616,
    g25431,II33257,g24909,II33260,g25436,g25437,g24627,g25438,II33265,g24925,
    II33268,g25443,g25444,g24641,g25445,g25449,g24660,II33278,g25088,g25454,
    II33282,g25096,g25458,II33286,g24426,g25462,II33289,g25106,g25463,II33293,
    g25008,g25467,II33297,g24430,g25471,II33300,g25112,g25472,II33304,g25004,
    g25476,II33307,g25011,g25479,II33312,g25014,g25484,II33316,g24434,g25488,
    II33321,g24442,g25493,II33324,g25009,g25496,II33327,g25017,g25499,II33330,
    g25019,g25502,II33335,g25010,g25507,II33338,g25021,g25510,II33343,g25024,
    g25515,II33347,g24438,g25519,II33352,g24443,g25524,II33355,g25012,g25527,
    II33358,g25028,g25530,II33361,g25013,g25533,II33364,g25029,g25536,II33368,
    g24444,g25540,II33371,g25015,g25543,II33374,g25031,g25546,II33377,g25033,
    g25549,II33382,g25016,g25554,II33385,g25035,g25557,II33390,g25038,g25562,
    II33396,g24447,g25573,II33399,g25018,g25576,II33402,g24448,g25579,II33405,
    g25020,g25582,II33408,g25040,g25585,II33411,g24491,g25588,II33415,g24449,
    g25590,II33418,g25022,g25593,II33421,g25043,g25596,II33424,g25023,g25599,
    II33427,g25044,g25602,II33431,g24450,g25606,II33434,g25025,g25609,II33437,
    g25046,g25612,II33440,g25048,g25615,II33445,g25026,g25620,II33448,g25050,
    g25623,g25630,g24478,II33457,g24451,g25634,II33460,g24452,g25637,II33463,
    g25030,g25640,II33466,g25053,g25643,II33469,g24498,g25646,II33472,g24499,
    g25647,II33476,g24453,g25652,II33479,g25032,g25655,II33482,g24454,g25658,
    II33485,g25034,g25661,II33488,g25054,g25664,II33491,g24501,g25667,II33495,
    g24455,g25669,II33498,g25036,g25672,II33501,g25057,g25675,II33504,g25037,
    g25678,II33507,g25058,g25681,II33511,g24456,g25685,II33514,g25039,g25688,
    II33517,g25060,g25691,II33520,g25062,g25694,g25698,II33526,g24457,g25700,
    II33529,g25041,g25703,II33532,g24507,g25706,II33535,g24508,g25707,II33539,
    g24458,g25711,II33542,g24459,g25714,II33545,g25045,g25717,II33548,g25064,
    g25720,II33551,g24510,g25723,II33554,g24511,g25724,II33558,g24460,g25729,
    II33561,g25047,g25732,II33564,g24461,g25735,II33567,g25049,g25738,II33570,
    g25065,g25741,II33573,g24513,g25744,II33577,g24462,g25746,II33580,g25051,
    g25749,II33583,g25068,g25752,II33586,g25052,g25755,II33589,g25069,g25758,
    II33593,g24445,g25762,II33596,g24446,g25763,II33600,g24463,g25767,II33603,
    g24519,g25770,g25771,II33608,g24464,g25773,II33611,g25055,g25776,II33614,
    g24521,g25779,II33617,g24522,g25780,II33621,g24465,g25784,II33624,g24466,
    g25787,II33627,g25059,g25790,II33630,g25071,g25793,II33633,g24524,g25796,
    II33636,g24525,g25797,II33640,g24467,g25802,II33643,g25061,g25805,II33646,
    g24468,g25808,II33649,g25063,g25811,II33652,g25072,g25814,II33655,g24527,
    g25817,II33659,g24469,g25821,II33662,g24532,g25824,g25825,II33667,g24470,
    g25827,II33670,g25066,g25830,II33673,g24534,g25833,II33676,g24535,g25834,
    II33680,g24471,g25838,II33683,g24472,g25841,II33686,g25070,g25844,II33689,
    g25074,g25847,II33692,g24537,g25850,II33695,g24538,g25851,II33700,g24474,
    g25856,II33703,g24545,g25859,g25860,II33708,g24475,g25862,II33711,g25073,
    g25865,II33714,g24547,g25868,II33717,g24548,g25869,II33723,g24477,g25877,
    II33726,g24557,g25880,II33732,g24473,g25886,II33737,g24476,g25891,g25895,
    g25899,g24928,g25903,g25907,g24940,g25911,g25915,g24951,g25919,g25923,
    g24963,g25937,g25939,g25942,g25945,g25952,II33790,g25976,II33798,g25982,
    II33801,II33804,II33807,II33810,II33813,II33816,II33819,II33822,II33825,
    II33828,II33831,II33834,II33837,II33840,II33843,II33846,II33849,II33852,
    II33855,II33858,II33861,II33864,II33867,II33870,II33873,II33876,II33879,
    II33882,II33885,II33888,II33891,II33894,II33897,II33900,II33903,II33906,
    II33909,II33912,II33915,II33918,II33954,g25343,g26056,II33961,g25357,
    g26063,II33968,g25372,g26070,II33974,g25389,g26076,II33984,g25932,g26086,
    II33990,g25870,g26092,II33995,g25935,g26102,II33999,g25490,II34002,g26105,
    II34009,g25882,g26114,II34012,g25938,g26118,II34017,g25887,g26121,II34020,
    g25940,g26125,II34026,g25892,g26131,II34029,g25520,II34032,g26136,II34041,
    g25566,II34044,g26150,II34051,g25204,g26159,II34056,g25206,g26164,II34059,
    g25207,g26165,II34063,g25209,g26167,II34068,g25211,g26172,II34071,g25212,
    g26173,II34074,g25213,g26174,II34077,g25954,g26175,II34080,g25539,g26178,
    II34083,g25214,g26181,II34086,g25215,g26182,II34091,g25217,g26187,g26189,
    II34096,g25218,g26190,II34099,g25219,g26191,II34102,g25220,g26192,II34105,
    g25221,g26193,II34108,g25222,g26194,II34111,g25223,g26195,II34114,g25958,
    g26196,II34118,g25605,g26202,II34121,g25224,g26205,II34124,g25225,g26206,
    II34128,g25227,g26208,g26209,II34132,g25228,g26210,II34135,g25229,g26211,
    II34140,g25230,g26214,II34143,g25231,g26215,II34146,g25232,g26216,II34150,
    g25233,g26220,II34153,g25234,g26221,II34156,g25235,g26222,II34159,g25964,
    g26223,II34162,g25684,g26226,II34165,g25236,g26229,II34168,g25237,g26230,
    II34172,g25239,g26232,g26237,II34180,g25240,g26238,II34183,g25241,g26239,
    II34189,g25242,g26245,II34192,g25243,g26246,II34195,g25244,g26247,II34198,
    g25245,g26248,II34201,g25246,g26249,II34204,g25247,g26250,II34207,g25969,
    g26251,II34210,g25761,g26254,II34220,g25248,g26264,g26275,II34230,g25249,
    g26276,II34233,g25250,g26277,II34238,g25251,g26280,II34241,g25252,g26281,
    II34244,g25253,g26282,II34254,g25185,g26294,II34266,g25255,g26308,g26313,
    II34274,g25256,g26314,II34277,g25257,g26315,II34296,g25189,g26341,II34306,
    g25259,g26349,II34313,g25265,g26354,II34316,g25191,g26355,II34321,g25928,
    g26358,II34327,g25260,g26364,II34343,g25194,g26385,II34353,g25927,g26393,
    II34358,g25262,g26398,II34363,g25930,g26401,II34369,g25263,g26407,II34385,
    g25197,g26428,II34388,g25200,g26429,II34392,g25266,g26433,II34395,g25929,
    g26434,II34400,g25267,g26439,II34405,g25933,g26442,II34411,g25268,g26448,
    II34421,g25203,g26461,II34425,g25270,g26465,II34428,g25931,g26466,II34433,
    g25271,g26471,II34438,g25936,g26474,II34444,g25272,g26480,g26481,g25764,
    II34449,g25205,g26485,II34453,g25279,g26489,II34456,g25934,g26490,II34461,
    g25280,g26495,II34464,g25199,g26496,g26497,g25818,II34469,g25210,g26501,
    II34473,g25288,g26505,II34476,g25201,g26506,II34479,g25202,g26507,g26508,
    g25312,g26512,g25853,g26516,g25320,g26520,g25874,g26521,g25331,g26525,
    g25340,g26533,g26538,g26539,g26540,g26542,g26543,g26544,g26546,II34505,
    g25450,g26548,g26549,g26550,g26551,g26552,g26554,g26555,g26556,g26558,
    g26561,g26562,g26563,g26564,g26565,g26566,g26567,g26568,g26570,g26571,
    g26572,g26574,II34535,g25451,g26576,g26577,g26578,g26579,g26580,g26581,
    g26582,g26584,g26585,g26586,g26587,g26588,g26589,g26590,g26591,g26593,
    g26594,g26595,g26597,g26598,g26599,g26600,g26601,g26602,g26603,g26604,
    g26605,g26606,g26608,g26609,g26610,g26611,g26612,g26613,g26614,g26615,
    g26617,II34579,g25452,g26618,g26619,g26620,g26621,g26622,g26623,g26624,
    g26625,g26626,g26627,g26628,g26629,g26631,g26632,g26633,g26634,g26635,
    g26636,g26637,g26638,g26639,g26640,g26641,g26642,g26643,g26644,g26645,
    g26646,g26647,g26648,g26649,g26650,g26651,g26652,g26653,g26654,g26656,
    g26657,g26658,g26662,II34641,II34644,II34647,II34650,II34653,II34656,
    II34659,II34662,II34665,II34668,II34671,II34674,II34677,II34680,II34683,
    II34686,II34689,II34692,II34695,II34698,II34701,II34704,II34707,II34710,
    II34713,II34716,II34719,II34722,II34725,II34728,II34731,II34734,II34737,
    II34740,II34743,II34746,II34749,II34752,II34755,II34758,II34761,II34764,
    II34767,II34770,II34773,II34776,II34779,II34782,II34785,II34788,II34791,
    II34794,II34797,II34800,II34803,II34806,II34809,II34812,II34815,II34818,
    II34821,II34824,II34827,II34830,II34833,II34836,II34839,II34842,II34845,
    II34848,II34851,II34854,II34857,II34860,II34863,II34866,II34872,g26217,
    g26757,II34879,g26240,g26762,II34901,g26295,g26782,II34909,g26265,g26788,
    II34916,g26793,II34921,g26796,II34946,g26534,g26819,II34957,g26541,g26828,
    II34961,g26545,g26830,II34964,g26547,g26831,II34967,g26553,g26832,II34971,
    g26557,g26834,II34974,g26168,g26835,II34977,g26559,g26836,II34980,g26458,
    g26837,II34983,g26569,g26840,II34986,g26160,g26841,II34990,g26573,g26843,
    II34993,g26575,g26844,II34997,g26482,g26846,II35000,g26336,g26849,II35003,
    g26592,g26850,II35007,g26596,g26852,II35011,g26304,g26854,II35014,g26498,
    g26855,II35017,g26616,g26858,II35028,g26513,g26861,II35031,g26529,g26864,
    II35049,g26530,g26868,II35053,g26655,g26872,II35064,g26531,g26875,II35067,
    g26659,g26876,II35072,g26661,g26881,II35076,g26532,g26883,II35079,g26664,
    g26884,II35083,g26665,g26886,II35087,g26667,g26890,II35092,g26669,g26895,
    II35095,g26670,g26896,II35099,g26672,g26900,II35106,g26675,g26909,II35109,
    g26676,g26910,II35116,g26025,g26921,g26922,g26283,g26935,g26327,g26944,
    g26374,g26950,g26417,II35136,g26660,g26953,g26954,II35141,g26666,g26956,
    g26957,II35146,g26671,g26959,g26960,II35153,g26677,g26964,II35172,g26272,
    g26983,g26987,g27010,g27036,g27064,II35254,g26048,g27075,II35283,g26031,
    g27102,II35297,g26199,g27114,II35301,g26037,g27116,II35313,g27126,II35319,
    g26183,g27132,g27133,g27134,g27135,g27136,g27137,g27138,g27139,g27140,
    g27141,g27142,g27143,II35334,g26106,g27145,g27146,g27148,II35341,g26120,
    g27150,g27151,g27153,II35347,g27154,g27155,II35351,g27156,II35355,g26130,
    g27158,g27159,II35360,g27161,g27162,II35364,g27163,g27164,II35369,g26144,
    g27166,g27167,II35373,g27168,II35376,g27171,g27172,g27173,II35383,g27176,
    g27177,II35389,g27180,II35394,g27183,II35399,g27186,II35404,II35407,
    II35410,II35413,II35416,II35419,II35422,II35425,II35428,II35431,II35434,
    II35437,II35440,II35443,II35446,II35449,II35452,II35455,II35458,II35461,
    II35464,II35467,II35470,II35473,II35476,II35479,II35482,II35485,II35488,
    II35491,II35494,II35497,II35500,II35503,II35506,II35509,II35512,II35515,
    II35518,II35521,II35524,II35527,II35530,II35533,II35536,II35539,II35542,
    II35545,II35548,II35551,II35554,g27349,II35667,g27120,g27353,II35673,
    g27123,g27357,II35678,g27129,g27360,II35681,g26869,g27361,II35686,g27131,
    g27366,II35689,g26878,g27367,II35695,g26887,g27373,II35698,g26897,g27376,
    II35708,g26974,II35711,g27381,g27383,g27384,II35723,g27385,g27386,II35727,
    g26902,g27387,II35731,g26892,g27391,II35737,g26915,g27397,II35741,g27118,
    g27401,II35744,g26906,g27404,II35750,g26928,g27410,II35756,g27117,g27416,
    II35759,g27121,g27419,II35762,g26918,g27422,II35768,g26941,g27428,II35772,
    g26772,g27432,II35777,g27119,g27437,II35780,g27124,g27440,II35783,g26931,
    g27443,g27449,II35791,g26779,g27451,II35796,g27122,g27456,II35799,g27130,
    g27459,II35803,g26803,g27463,g27465,II35809,g26785,g27467,II35814,g27125,
    g27472,II35817,g27475,II35821,g26804,g27479,II35824,g26805,g27480,II35829,
    g26806,g27483,g27484,II35834,g26792,g27486,II35837,g26911,g27489,II35841,
    g26807,g27493,II35844,g26808,g27494,II35849,g26776,g27497,II35852,g27498,
    II35856,g26809,g27502,II35859,g26810,g27503,II35863,g26811,g27505,g27506,
    II35868,g26812,g27508,II35872,g26925,g27510,II35876,g26813,g27514,II35879,
    g26814,g27515,II35883,g26781,g27517,II35886,g27518,II35890,g26815,g27522,
    II35893,g26816,g27523,II35897,g26817,g27525,II35900,g26786,g27526,II35915,
    g26818,g27533,II35919,g26938,g27535,II35923,g26820,g27539,II35926,g26821,
    g27540,II35930,g26789,g27542,II35933,g27543,II35937,g26822,g27547,II35940,
    g26823,g27548,II35953,g26824,g27553,II35957,g26947,g27555,II35961,g26825,
    g27559,II35964,g26826,g27560,II35968,g26795,g27562,II35983,g26827,g27569,
    II36008,g26798,g27586,g27589,g27590,g27144,g27595,g27149,g27599,g27147,
    g27604,g27157,g27608,g27152,g27613,g27165,g27617,g27160,g27622,g27174,
    II36032,g27113,g27632,II36042,g27662,II36046,g27667,II36052,g27674,II36060,
    II36063,II36066,II36069,II36072,II36075,II36078,II36081,II36084,II36087,
    II36090,II36093,II36096,II36099,II36102,II36105,II36108,II36111,II36114,
    II36117,II36120,II36123,II36126,II36129,II36132,II36135,II36138,II36141,
    II36144,II36147,II36150,II36153,II36156,II36159,II36162,g27748,II36213,
    g27571,g27776,II36217,g27580,g27780,II36221,g27784,II36224,g27785,II36227,
    g27594,g27786,II36230,g27583,g27787,II36234,g27791,II36237,g27792,II36240,
    g27603,g27793,II36243,g27587,g27794,II36246,g27797,II36250,g27612,g27799,
    II36253,g27800,II36264,g27621,g27805,II36267,g27395,g27806,II36280,g27390,
    g27817,II36283,g27408,g27820,II36296,g27626,g27831,II36307,g27400,g27839,
    II36311,g27426,g27843,II36321,g27627,g27847,II36327,g27413,g27858,II36330,
    g27447,g27861,II36337,g27628,g27872,II36341,g27431,g27879,II36347,g27630,
    g27889,II36354,g27903,II36358,g27672,g27905,II36362,g27907,II36367,g27678,
    g27910,II36371,g27912,II36379,g27682,g27918,II36382,g27563,g27919,II36390,
    g27243,g27927,II36393,g27572,g27928,II36397,g27574,g27932,II36404,g27450,
    g27939,II36407,g27581,g27942,II36411,g27582,g27946,II36417,g27462,g27952,
    II36420,g27253,g27955,II36423,g27466,g27956,II36426,g27584,g27959,II36432,
    g27585,g27965,g27969,II36438,g27255,g27971,II36441,g27256,g27972,II36444,
    g27482,g27973,II36447,g27257,g27976,II36450,g27485,g27977,II36454,g27588,
    g27981,II36459,g27258,g27986,II36462,g27259,g27987,II36465,g27260,g27988,
    II36468,g27261,g27989,g27990,II36473,g27262,g27992,II36476,g27263,g27993,
    II36479,g27504,g27994,II36483,g27264,g27998,II36486,g27507,g27999,II36490,
    g27265,g28003,II36493,g27266,g28004,II36496,g27267,g28005,II36499,g27268,
    g28006,II36502,g27269,g28007,II36507,g27270,g28010,II36510,g27271,g28011,
    II36513,g27272,g28012,II36516,g27273,g28013,g28014,II36521,g27274,g28016,
    II36524,g27275,g28017,II36527,g27524,g28018,II36530,g27276,g28021,II36533,
    g27277,g28022,II36536,g27278,g28023,II36539,g27279,g28024,II36542,g27280,
    g28025,II36545,g27281,g28026,II36551,g27282,g28030,II36554,g27283,g28031,
    II36557,g27284,g28032,II36560,g27285,g28033,II36563,g27286,g28034,II36568,
    g27287,g28037,II36571,g27288,g28038,II36574,g27289,g28039,II36577,g27290,
    g28040,g28041,II36582,g27291,g28043,II36585,g27292,g28044,II36588,g27293,
    g28045,II36598,g27294,g28047,II36601,g27295,g28048,II36604,g27296,g28049,
    II36609,g27297,g28052,II36612,g27298,g28053,II36615,g27299,g28054,II36618,
    g27300,g28055,II36621,g27301,g28056,II36627,g27302,g28060,II36630,g27303,
    g28061,II36633,g27304,g28062,II36636,g27305,g28063,II36639,g27306,g28064,
    II36644,g27307,g28067,II36647,g27308,g28068,II36650,g27309,g28069,II36653,
    g27310,g28070,II36656,g27311,g28071,II36659,g27312,g28072,II36663,g27313,
    g28074,II36673,g27314,g28076,II36676,g27315,g28077,II36679,g27316,g28078,
    II36684,g27317,g28081,II36687,g27318,g28082,II36690,g27319,g28083,II36693,
    g27320,g28084,II36696,g27321,g28085,II36702,g27322,g28089,II36705,g27323,
    g28090,II36708,g27324,g28091,II36711,g27325,g28092,II36714,g27326,g28093,
    II36718,g27327,g28095,II36721,g27328,g28096,II36724,g27329,g28097,II36728,
    g27330,g28099,II36738,g27331,g28101,II36741,g27332,g28102,II36744,g27333,
    g28103,II36749,g27334,g28106,II36752,g27335,g28107,II36755,g27336,g28108,
    II36758,g27337,g28109,II36761,g27338,g28110,II36766,g27339,g28113,II36769,
    g27340,g28114,II36772,g27341,g28115,II36776,g27342,g28117,II36786,g27343,
    g28119,II36789,g27344,g28120,II36792,g27345,g28121,II36797,g27346,g28124,
    II36800,g27347,g28125,II36803,g27348,g28126,g28128,g27528,II36808,g27354,
    g28132,g28133,g27550,g28137,g27566,g28141,g27576,g28149,g28150,g28151,
    g28152,g28153,g28154,g28155,g28156,g28158,g28159,g28160,g28161,g28162,
    g28163,g28164,g28165,g28166,g28167,g28168,g28169,g28170,g28172,g28173,
    g28174,g28175,g28177,g28178,II36848,g28179,g28186,g28187,g28190,II36860,
    g28194,II36864,g28200,II36867,II36870,II36873,II36876,II36879,II36882,
    II36885,II36888,II36891,II36894,II36897,II36900,II36903,II36906,II36909,
    II36912,II36915,II36918,II36921,II36924,II36927,II36930,II36933,II36936,
    II36939,II36942,II36945,II36948,II36951,II36954,II36957,II36960,II36963,
    II36966,II36969,II36972,II36975,II36978,II36981,II36984,II36987,II36990,
    II36993,II36996,II36999,II37002,II37005,II37008,II37011,II37014,II37017,
    II37020,II37023,II37026,II37029,II37032,II37035,II37038,II37041,II37044,
    II37047,II37050,II37053,II37056,II37059,II37062,II37065,II37068,II37071,
    II37074,II37077,II37080,II37083,II37086,II37089,II37092,II37095,II37098,
    II37101,II37104,II37107,II37110,II37113,II37116,II37119,II37122,II37125,
    II37128,II37131,II37134,II37137,II37140,II37143,II37146,II37149,II37152,
    II37155,II37158,II37161,II37164,II37167,II37170,II37173,II37176,II37179,
    II37182,II37185,II37188,II37191,II37194,II37197,II37200,II37203,II37228,
    g28341,II37232,g28343,II37238,g28347,II37252,g28359,II37260,g28365,II37266,
    g28369,II37269,g28145,g28370,II37273,g28372,II37277,g28146,g28374,II37280,
    g28375,II37284,g28147,g28377,II37291,g28148,g28382,II37319,g28390,II37330,
    g28393,II37334,g28395,g28419,II37379,g28199,g28432,II37386,g28437,II37394,
    g27718,g28443,II37400,g28447,II37410,g27722,g28455,II37415,g28458,II37426,
    g27724,g28467,g28483,g28491,g28496,II37459,g27759,g28498,g28500,II37467,
    g27760,g28524,II37471,g27761,g28526,II37474,g27762,g28527,II37481,g27763,
    g28552,II37484,g27764,g28553,g28554,II37488,g27765,g28555,II37494,g27766,
    g28579,II37497,g27767,g28580,g28581,g28582,II37502,g27768,g28583,II37508,
    g27769,g28607,g28608,g28609,g28610,II37514,g27771,g28611,g28612,g28046,
    g28616,g28617,g28618,g28619,g28075,g28623,g28624,g28625,g28100,g28629,
    g28630,g28118,g28638,g28639,g28640,g28641,g28642,g28643,g28644,g28645,
    g28646,g28647,g28648,g28649,g28650,g28651,g28652,g28653,g28655,II37566,
    II37569,II37572,II37575,II37578,II37581,II37584,II37587,II37590,II37593,
    II37596,II37599,II37602,II37605,II37608,II37611,II37614,II37617,II37620,
    II37623,II37626,II37629,II37632,II37635,II37638,II37641,II37644,II37647,
    II37650,II37653,II37656,II37659,II37662,II37665,g28720,g28495,g28721,
    g28490,g28723,g28528,g28725,g28499,g28727,g28489,g28730,g28470,g28734,
    g28525,g28740,g28488,II37702,g28512,g28741,II37712,g28751,II37716,g28540,
    g28755,II37725,g28764,II37729,g28567,g28768,II37736,g28775,II37740,g28595,
    g28779,II37746,g28785,II37752,g28791,II37757,g28796,II37760,g28799,II37765,
    g28804,II37768,g28807,II37771,g28810,II37775,g28814,II37778,g28817,II37781,
    g28820,II37784,g28823,II37787,g28826,II37790,g28829,II37793,g28832,II37796,
    g28634,g28833,II37800,g28635,g28835,II37804,g28636,g28837,II37808,g28637,
    g28839,g28855,g28409,g28859,g28413,g28863,g28417,g28867,g28418,II37842,
    g28501,g28871,II37846,g28877,II37851,g28668,g28882,II37854,g28529,g28883,
    II37858,g28889,II37863,g28894,II37868,g28321,g28899,II37871,g28556,g28900,
    II37875,g28906,II37880,g28911,II37885,g28916,II37891,g28325,g28924,II37894,
    g28584,g28925,II37897,g28928,II37901,g28932,II37906,g28937,II37912,g28945,
    II37917,g28328,g28950,II37920,g28951,II37924,g28955,II37928,g28959,II37934,
    g28967,II37939,g28972,II37942,g28975,II37946,g28979,II37950,g28983,II37956,
    g28993,II37961,g28998,II37965,g29002,II37968,g29005,II37973,g29010,II37978,
    g29019,II37982,g29023,II37986,g29027,II37991,g29032,II37994,g29035,II37999,
    g29042,II38003,g29046,II38007,g29050,II38011,g29054,II38014,g29057,II38018,
    g28342,g29061,II38024,g29065,II38028,g29069,II38032,g28344,g29073,II38035,
    g28345,g29074,II38038,g28346,g29075,II38042,g29077,II38046,g28348,g29081,
    II38049,g28349,g29082,II38053,g28350,g29084,II38056,g28351,g29085,II38059,
    g28352,g29086,II38064,g28353,g29089,II38068,g28354,g29091,II38071,g28355,
    g29092,II38074,g28356,g29093,II38077,g28357,g29094,II38080,g28358,g29095,
    II38085,g28360,g29098,II38088,g28361,g29099,II38091,g28362,g29100,II38094,
    g28363,g29101,II38097,g28364,g29102,II38101,g28366,g29104,II38104,g28367,
    g29105,II38107,g28368,g29106,II38111,g28371,g29108,II38119,g28420,g29117,
    II38122,g28421,g29118,II38125,g28425,g29119,II38128,g29120,II38136,II38139,
    II38142,II38145,II38148,II38151,II38154,II38157,II38160,II38163,II38166,
    II38169,II38172,II38175,II38178,II38181,II38184,II38187,II38190,II38193,
    II38196,II38199,II38202,II38205,II38208,II38211,II38214,II38217,II38220,
    II38223,II38226,II38229,II38232,II38235,II38238,II38241,II38245,g28920,
    g29168,II38250,g28941,g29171,II38258,g28963,g29177,II38272,g29013,g29189,
    II38275,g28987,g29190,II38278,g29191,g29192,g28954,II38282,g29193,II38321,
    g29113,g29230,II38330,g29237,II38339,g29244,II38342,g28886,g29245,II38345,
    g29109,g29246,II38348,g28874,g29247,II38352,g29110,g29249,II38355,g29039,
    g29250,II38360,g29111,g29253,II38363,g29016,g29254,II38369,g29112,g29258,
    g29266,II38386,g29267,g29268,g29269,II38391,g29270,g29271,g29272,II38396,
    g29273,g29274,g29275,II38401,g29276,g29277,II38405,g29278,II38408,g29279,
    g29280,II38412,g29281,g29282,g29283,g29285,g29286,g29287,II38421,g29288,
    g29290,g29291,g29292,II38428,g28732,g29293,g29295,g29296,II38434,g28735,
    g29297,II38437,g28736,g29298,II38440,g28738,g29299,g29301,II38447,g28744,
    g29304,II38450,g28745,g29305,II38453,g28746,g29306,II38456,g28747,g29307,
    II38459,g28749,g29308,II38462,g29309,II38466,g28754,g29311,II38471,g28758,
    g29314,II38474,g28759,g29315,II38477,g28760,g29316,II38480,g28761,g29317,
    II38483,g28990,g29318,II38486,g28763,g29319,II38491,g28767,g29322,II38496,
    g28771,g29325,II38499,g28772,g29326,II38502,g28773,g29327,II38505,g28774,
    g29328,II38510,g28778,g29331,II38515,g28782,g29334,II38518,g28783,g29335,
    II38524,g28788,g29339,II38536,g29349,II38539,g29350,g29356,g29358,II38548,
    g28903,g29359,g29360,g29361,g29362,g29363,g29364,g29365,g29366,g29367,
    g29368,g29369,g29370,g29371,g29372,g29373,g29374,g29375,g29376,g29377,
    g29378,g29379,g29380,g29381,g29382,g29383,g29384,g29385,g29386,g29387,
    g29388,g29389,g29390,g29391,g29392,g29393,g29394,g29395,g29396,g29397,
    g29398,II38591,g29400,II38594,g29401,g29402,II38599,g29404,II38602,g29405,
    II38606,g29407,II38609,g29408,II38613,g29410,II38617,g29412,II38620,
    II38623,II38626,II38629,II38632,II38635,II38638,II38641,II38644,II38647,
    II38650,II38653,II38656,II38659,II38662,II38665,II38668,II38671,II38674,
    II38677,II38680,II38683,II38686,II38689,II38692,II38695,II38698,II38701,
    II38704,II38707,II38710,II38713,II38716,II38719,II38722,II38725,II38728,
    II38731,II38734,II38737,II38740,II38743,II38746,II38749,II38752,II38755,
    II38758,II38761,II38764,II38767,II38770,g29491,II38801,g29495,II38804,
    g29353,g29496,II38807,g29497,II38817,g29354,g29499,II38827,g29355,g29501,
    II38838,g29357,g29504,II38848,g29167,g29506,II38851,g29169,g29507,II38854,
    g29170,g29508,II38857,g29172,g29509,II38860,g29173,g29510,II38863,g29178,
    g29511,II38866,g29179,g29512,II38869,g29181,g29513,II38872,g29182,g29514,
    II38875,g29184,g29515,II38878,g29185,g29516,II38881,g29187,g29517,II38885,
    g29519,II38898,g29194,g29530,II38905,g29197,g29535,II38909,g29198,g29537,
    II38916,g29201,g29542,II38920,g29204,g29544,II38924,g29205,g29546,II38931,
    g29209,g29551,II38936,g29212,g29554,II38940,g29213,g29556,II38947,g29218,
    g29561,II38951,g29221,g29563,II38958,g29226,g29568,II38975,g29348,g29583,
    II38999,II39002,II39005,II39008,II39011,II39014,II39017,II39020,II39023,
    II39026,II39029,II39032,II39035,II39038,II39041,II39044,II39047,II39050,
    II39053,II39056,II39059,II39062,II39065,II39068,II39071,II39074,II39077,
    II39080,II39083,II39086,II39089,g29658,g29574,g29659,g29571,g29660,g29578,
    g29661,g29576,g29662,g29570,g29664,g29552,g29666,g29577,g29668,g29569,
    g29673,II39121,g29579,g29689,II39124,g29606,g29690,II39127,g29608,g29691,
    II39130,g29580,g29692,II39133,g29609,g29693,II39136,g29611,g29694,II39139,
    g29612,g29695,II39142,g29581,g29696,II39145,g29613,g29697,II39148,g29616,
    g29698,II39151,g29617,g29699,II39154,g29582,g29700,II39157,g29618,g29701,
    II39160,g29620,g29702,II39164,g29621,g29704,II39168,g29623,g29708,g29716,
    g29498,g29724,g29500,g29726,g29503,g29739,g29505,II39234,II39237,II39240,
    II39243,II39246,II39249,II39252,II39255,II39258,II39261,II39264,II39267,
    II39270,II39273,II39276,II39279,g29823,g29663,g29829,g29665,g29835,g29667,
    g29840,g29669,g29844,g29670,g29848,g29761,g29849,g29671,g29853,g29672,
    g29857,g29676,g29861,g29677,g29865,g29678,g29869,g29679,g29873,g29680,
    g29877,g29681,g29881,g29682,g29885,g29683,g29889,g29684,g29893,g29685,
    g29897,g29686,g29901,g29687,g29905,g29688,II39398,g29932,II39401,g29933,
    II39404,g29934,II39407,g29935,II39411,g29937,II39414,g29938,II39418,g29940,
    II39423,g29943,II39454,II39457,II39460,II39463,II39466,II39469,II39472,
    II39475,g30036,g29912,g30040,g29914,g30044,g29916,g30048,g29920,II39550,
    g30052,II39573,g29936,g30076,II39577,g29939,g30078,II39585,g29941,g30084,
    II39622,II39625,II39628,II39631,II39635,g30055,g30124,II39638,g30056,
    g30125,II39641,g30057,g30126,II39647,g30058,g30130,g30134,g30010,g30139,
    g30011,g30143,g30012,g30147,g30013,g30151,g30014,g30155,g30015,g30159,
    g30016,g30163,g30017,g30167,g30018,g30171,g30019,g30175,g30020,g30179,
    g30021,g30183,g30022,g30187,g30023,g30191,g30024,g30195,g30025,g30199,
    g30026,g30203,g30027,g30207,g30028,g30211,g30029,II39674,g30072,g30215,
    g30229,g30030,g30233,g30031,g30237,g30032,g30241,g30033,II39761,g30306,
    II39764,g30060,g30307,II39767,g30061,g30308,II39770,g30063,g30309,II39773,
    g30064,g30310,II39776,g30066,g30311,II39779,g30053,g30312,II39782,g30054,
    g30313,II39785,II39788,II39791,II39794,II39797,II39800,II39803,II39806,
    II39809,II39812,II39815,II39818,II39821,g30267,g30326,II39825,g30268,
    g30328,II39828,g30269,g30329,II39832,g30270,g30331,II39835,g30271,g30332,
    II39840,g30272,g30335,II39843,g30273,g30336,II39848,g30274,g30339,II39853,
    g30275,g30342,II39856,g30276,g30343,II39859,g30277,g30344,II39863,g30278,
    g30346,II39866,g30279,g30347,II39870,g30280,g30349,II39873,g30281,g30350,
    II39878,g30282,g30353,II39881,g30283,g30354,II39886,g30284,g30357,II39889,
    g30285,g30358,II39892,g30286,g30359,II39895,g30287,g30360,II39899,g30288,
    g30362,II39902,g30289,g30363,II39906,g30290,g30365,II39909,g30291,g30366,
    II39913,g30292,g30368,II39916,g30293,g30369,II39919,g30294,g30370,II39922,
    g30295,g30371,II39926,g30296,g30373,II39930,g30297,g30375,II39933,g30298,
    g30376,II39936,g30299,g30377,II39939,g30300,g30378,II39942,g30301,g30379,
    II39945,g30302,g30380,II39948,g30303,g30381,II39951,g30304,g30382,g30383,
    II39976,g30245,g30408,II39982,g30305,g30412,II39985,g30246,g30435,II39991,
    g30247,g30439,II39997,g30248,g30443,II40002,g30249,g30446,II40008,g30250,
    g30450,II40016,g30251,g30456,II40021,g30252,g30459,II40027,g30253,g30463,
    II40032,g30254,g30466,II40039,g30255,g30471,II40044,g30256,g30474,II40051,
    g30257,g30479,II40054,g30258,g30480,II40059,g30259,g30483,II40066,g30260,
    g30488,II40071,g30261,g30491,II40075,g30262,g30493,II40078,g30263,g30494,
    II40083,g30264,g30497,II40086,g30265,g30498,II40091,g30266,g30501,II40098,
    II40101,II40104,II40107,II40110,II40113,II40116,II40119,II40122,II40125,
    II40128,II40131,II40134,II40137,II40140,II40143,II40146,II40149,II40152,
    II40155,II40158,II40161,II40164,II40167,II40170,II40173,II40176,II40179,
    II40182,II40185,II40188,II40191,II40194,II40197,II40200,II40203,II40206,
    II40209,II40212,II40215,II40218,II40221,II40224,II40227,II40230,II40233,
    II40236,II40239,II40242,II40245,II40248,II40251,II40254,II40257,II40260,
    II40263,II40266,II40269,II40272,II40275,g30567,g30403,g30568,g30402,g30569,
    g30406,g30570,g30404,g30571,g30401,g30572,g30399,g30573,g30405,g30574,
    g30400,g30575,II40288,g30455,g30578,II40291,g30468,g30579,II40294,g30470,
    g30580,II40297,g30482,g30581,II40300,g30485,g30582,II40303,g30487,g30583,
    II40307,g30500,g30585,II40310,g30503,g30586,II40313,g30505,g30587,II40317,
    g30338,g30591,II40320,g30341,g30592,II40326,g30356,g30600,II40420,II40423,
    II40426,II40429,II40432,II40435,II40438,II40441,II40444,II40447,II40450,
    II40453,II40456,g30668,g30722,II40459,g30669,g30723,II40462,g30670,g30724,
    II40465,g30671,g30725,II40468,g30672,g30726,II40471,g30673,g30727,II40475,
    g30674,g30729,II40478,g30675,g30730,II40481,g30676,g30731,II40484,g30677,
    g30732,II40487,g30678,g30733,II40490,g30679,g30734,II40495,g30680,g30737,
    II40498,g30681,g30738,II40501,g30682,g30739,II40504,g30683,g30740,II40507,
    g30684,g30741,II40510,g30686,g30742,II40515,g30687,g30745,II40518,g30688,
    g30746,II40521,g30689,g30747,II40524,g30690,g30748,II40527,g30691,g30749,
    II40531,g30692,g30751,II40534,g30693,g30752,II40537,g30694,g30753,II40542,
    g30695,g30756,g30765,g30685,II40555,g30699,g30767,II40565,g30700,g30769,
    II40568,g30701,g30770,II40578,g30702,g30772,II40581,g30703,g30773,II40584,
    g30704,g30774,II40594,g30705,g30776,II40597,g30706,g30777,II40600,g30707,
    g30778,II40611,g30708,g30781,II40614,g30709,g30782,II40618,g30566,g30784,
    II40634,g30792,II40637,g30793,II40640,g30794,II40643,g30795,II40647,g30797,
    II40651,g30799,II40654,g30800,II40658,g30802,II40661,g30635,g30803,II40664,
    g30636,g30804,II40667,g30637,g30805,II40670,g30638,g30806,II40673,g30639,
    g30807,II40676,g30640,g30808,II40679,g30641,g30809,II40682,g30642,g30810,
    II40685,g30643,g30811,II40688,g30644,g30812,II40691,g30645,g30813,II40694,
    g30646,g30814,II40697,g30647,g30815,II40700,g30648,g30816,II40703,g30649,
    g30817,II40706,g30650,g30818,II40709,g30651,g30819,II40712,g30652,g30820,
    II40715,g30653,g30821,II40718,g30654,g30822,II40721,g30655,g30823,II40724,
    g30656,g30824,II40727,g30657,g30825,II40730,g30658,g30826,II40733,g30659,
    g30827,II40736,g30660,g30828,II40739,g30661,g30829,II40742,g30662,g30830,
    II40745,g30663,g30831,II40748,g30664,g30832,II40751,g30665,g30833,II40754,
    g30666,g30834,II40757,g30667,g30835,II40760,II40763,II40766,II40769,
    II40772,II40775,II40778,II40781,II40784,II40787,II40790,II40793,II40796,
    II40799,II40802,II40805,II40808,II40811,II40814,II40817,II40820,II40823,
    II40826,II40829,II40832,II40835,II40838,II40841,II40844,II40847,II40850,
    II40853,II40856,II40859,II40862,II40865,II40868,II40871,II40874,II40877,
    II40880,II40883,II40886,II40889,II40892,II40895,II40898,II40901,II40904,
    II40907,II40910,II40913,II40916,II40919,II40922,II40925,II40928,II40931,
    II40934,II40937,II40940,II40943,II40946,II40949,II40952,II40955,II40958,
    II40961,II40964,II40967,II40970,II40973,II40976,II40979,II40982,II40985,
    II40988,II40991,II40994,II40997,II41024,g30928,II41035,g30796,g30937,
    II41038,g30798,g30938,II41041,g30801,g30939,II41044,II41047,II41050,
    II41053,g30962,g30958,g30963,g30957,g30964,g30961,g30965,g30959,g30966,
    g30956,g30967,g30954,g30968,g30960,g30969,g30955,g30971,g30970,II41090,
    g30972,II41093,g30973,II41096,g30974,II41099,g30975,II41102,g30976,II41105,
    g30977,II41108,g30978,II41111,g30979,II41114,II41117,II41120,II41123,
    II41126,II41129,II41132,II41135,II41138,g30988,II41141,g5630,g5649,g5650,
    g5658,g5676,g5677,g5678,g5687,g5688,g5696,g5709,g5710,g5711,g5728,g5729,
    g5730,g5739,g5740,g5748,g5757,g5758,g5767,g5768,g5769,g5786,g5787,g5788,
    g5797,g5798,g5807,g5816,g5817,g5826,g5827,g5828,g5845,g5846,g5847,g5863,
    g5872,g5873,g5882,g5883,g5884,g5910,g5919,g5920,g5949,g8327,g8328,g8329,
    g8339,g8340,g8350,g8385,g8386,g8387,g8394,g8395,g8396,g8406,g8407,g8417,
    g8431,g8432,g8433,g8437,g8438,g8439,g8446,g8447,g8448,g8458,g8459,g8463,
    g8464,g8465,g8466,g8467,g8468,g8472,g8473,g8474,g8481,g8482,g8483,g8484,
    g8485,g8486,g8487,g8488,g8489,g8490,g8491,g8492,g8493,g8497,g8498,g8499,
    g8500,g8501,g8502,g8503,g8504,g8505,g8506,g8507,g8508,g8509,g8510,g8511,
    g8512,g8513,g8515,g8516,g8517,g8518,g8519,g8520,g8521,g8522,g8523,g8524,
    g8525,g8526,g8527,g8528,g8529,g8531,g8532,g8534,g8535,g8536,g8537,g8538,
    g8539,g8540,g8541,g8542,g8543,g8544,g8545,g8546,g8548,g8549,g8551,g8552,
    g8553,g8554,g8555,g8556,g8557,g8558,g8559,g8561,g8562,g8564,g8565,g8566,
    g8567,g8570,g8572,g8573,g8576,g8601,g8612,g8613,g8621,g8625,g8626,g8631,
    g8635,g8636,g8650,g8654,g8666,g8676,g8687,g8688,g8703,g8704,g8705,g8706,
    g8717,g8722,g8723,g8724,g8725,g8751,g8755,g8760,g8761,g8762,g8774,g8778,
    g8783,g8784,g8797,g8801,g8816,g8841,g8842,g8861,g8868,g8869,g8892,g8899,
    g8906,g8907,g8932,g8939,g8946,g8947,g8972,g8979,g9004,g9009,g9026,g9033,
    g9034,g9047,g9048,g9049,g9056,g9057,g9061,g9062,g9063,g9064,g9065,g9066,
    g9073,g9074,g9075,g9076,g9077,g9078,g9079,g9080,g9081,g9082,g9083,g9090,
    g9091,g9092,g9093,g9094,g9095,g9096,g9097,g9098,g9099,g9100,g9101,g9102,
    g9103,g9104,g9105,g9106,g9107,g9108,g9109,g9110,g9111,g9112,g9113,g9114,
    g9115,g9116,g9117,g9118,g9119,g9120,g9121,g9122,g9123,g9124,g9125,g9126,
    g9127,g9131,g9132,g9133,g9137,g9138,g9139,g9143,g9145,g9241,g9301,g9302,
    g9319,g9364,g9365,g9366,g9367,g9382,g9383,g9400,g9438,g9439,g9440,g9441,
    g9442,g9461,g9462,g9463,g9464,g9479,g9480,g9497,g9518,g9519,g9520,g9521,
    g9522,g9523,g9534,g9580,g9581,g9582,g9583,g9584,g9603,g9604,g9605,g9606,
    g9621,g9622,g9630,g9631,g9632,g9633,g9634,g9635,II16735,II16736,g9636,
    g9639,g9647,g9648,g9660,g9661,g9662,g9663,g9664,g9665,g9676,g9722,g9723,
    g9724,g9725,g9726,g9745,g9746,g9747,g9748,g9759,g9760,g9761,g9762,g9763,
    g9764,g9765,g9766,g9773,g9774,g9775,g9776,g9777,g9778,g9779,g9780,g9781,
    II16826,II16827,g9782,g9785,g9793,g9794,g9806,g9807,g9808,g9809,g9810,
    g9811,g9822,g9868,g9869,g9870,g9871,g9872,g9887,g9888,g9889,g9890,g9891,
    g9892,g9893,g9894,g9901,g9902,g9903,g9904,g9905,g9906,g9907,g9908,g9909,
    g9910,g9911,g9912,g9919,g9920,g9921,g9922,g9923,g9924,g9925,g9926,g9927,
    II16930,II16931,g9928,g9931,g9939,g9940,g9952,g9953,g9954,g9955,g9956,
    g9957,g9968,g10007,g10008,g10009,g10010,g10011,g10012,g10013,g10014,g10024,
    g10035,g10036,g10037,g10041,g10042,g10043,g10044,g10045,g10046,g10047,
    g10048,g10055,g10056,g10057,g10058,g10059,g10060,g10061,g10062,g10063,
    g10064,g10065,g10066,g10073,g10074,g10075,g10076,g10077,g10078,g10079,
    g10080,g10081,II17042,II17043,g10082,g10085,g10093,g10094,g10101,g10102,
    g10103,g10104,g10105,g10106,g10107,g10108,g10112,g10113,g10114,g10115,
    g10116,g10117,g10118,g10119,g10120,g10121,g10122,g10123,g10133,g10144,
    g10145,g10146,g10150,g10151,g10152,g10153,g10154,g10155,g10156,g10157,
    g10164,g10165,g10166,g10167,g10168,g10169,g10170,g10171,g10172,g10173,
    g10174,g10175,g10182,g10183,g10184,II17156,g10186,g10192,g10193,g10194,
    g10195,g10196,g10197,g10198,g10199,g10200,g10201,g10202,g10203,g10204,
    g10205,g10206,g10207,g10208,g10209,g10210,g10211,g10212,g10213,g10217,
    g10218,g10219,g10220,g10221,g10222,g10223,g10224,g10225,g10226,g10227,
    g10228,g10238,g10249,g10250,g10251,g10255,g10256,g10257,g10258,g10259,
    g10260,g10261,g10262,g10269,g10270,g10271,g10272,g10279,g10280,g10281,
    g10282,g10283,g10284,g10285,g10286,g10287,g10288,g10289,g10290,g10291,
    g10292,g10293,g10294,g10295,g10296,g10297,g10298,g10299,g10300,g10301,
    g10302,g10303,g10304,g10305,g10306,g10307,g10308,g10309,g10310,g10311,
    g10312,g10313,g10314,g10315,g10319,g10320,g10321,g10322,g10323,g10324,
    g10325,g10326,g10327,g10328,g10329,g10330,g10340,g10351,g10352,g10353,
    g10360,g10361,g10362,g10363,g10364,g10365,g10366,g10367,g10368,g10369,
    g10370,g10371,g10372,g10373,g10374,g10375,g10376,g10377,g10378,g10379,
    g10380,g10381,g10382,g10383,g10384,g10385,g10386,g10387,g10388,g10389,
    g10390,g10391,g10392,g10393,g10394,g10395,g10396,g10397,g10398,g10399,
    g10400,g10401,g10402,g10403,g10404,g10405,g10406,g10407,g10408,g10412,
    g10413,g10414,g10415,g10422,g10423,g10430,g10431,g10432,g10433,g10434,
    g10435,g10436,g10437,g10438,g10439,g10440,g10441,g10442,g10443,g10444,
    g10445,g10446,g10447,g10448,g10449,g10450,g10451,g10452,g10453,g10454,
    g10455,g10456,g10457,g10458,g10459,g10460,g10461,g10462,g10463,g10464,
    g10465,g10466,g10467,g10468,g10469,g10470,g10471,g10472,g10473,g10474,
    g10475,g10476,g10477,g10478,g10479,II17429,g10485,g10492,g10493,g10494,
    g10495,g10496,g10497,g10498,g10499,g10506,g10507,g10508,g10509,g10510,
    g10511,g10512,g10513,g10514,g10515,g10516,g10517,g10518,g10519,g10520,
    g10521,g10522,g10523,g10524,g10525,g10526,g10527,g10528,g10529,g10530,
    g10531,g10532,g10533,g10534,g10535,g10536,g10537,g10538,g10539,g10540,
    g10541,g10548,g10555,g10556,g10557,g10558,g10559,g10566,g10567,g10568,
    g10569,g10570,g10571,g10572,g10573,g10580,g10581,g10582,g10583,g10584,
    g10585,g10586,g10587,g10588,g10589,g10590,g10591,g10592,g10593,g10594,
    g10595,g10596,g10597,g10598,g10599,g10600,g10604,g10605,g10612,g10613,
    g10614,g10615,g10616,g10623,g10624,g10625,g10626,g10627,g10628,g10629,
    g10630,g10637,g10638,g10639,g10640,g10641,g10642,g10643,g10644,g10645,
    g10650,g10651,g10652,g10659,g10660,g10661,g10662,g10663,g10670,g10671,
    g10672,g10673,g10674,g10675,g10678,g10680,g10681,g10682,g10689,g10690,
    g10691,g10692,g10693,g10704,g10707,g10709,g10710,II17599,g10724,g10727,
    g10729,g10745,g10748,g10764,g11347,g11420,g11421,g11431,g11607,g11612,
    g11637,g11771,g11788,g11805,g11814,g11816,g11838,g11847,g11851,g11880,
    g11885,g11922,g11926,g11966,g11967,g12012,g12069,g12070,g12128,g12129,
    g12186,g12273,g12274,g12307,g12330,g12331,g12353,g12376,g12419,g12429,
    g12477,g12494,g12514,g12531,g12650,II19937,II19938,g12876,g12908,II19971,
    II19972,g12916,g12938,II19996,II19997,g12945,g12966,II20021,II20022,g12974,
    g12989,g12990,g13000,g13009,g13010,g13023,g13031,g13032,g13042,II20100,
    g13056,II20131,II20132,g13247,g13266,g13270,g13289,g13291,g13295,g13316,
    g13320,g13322,g13326,g13335,g13340,g13343,g13345,g13355,g13360,g13365,
    g13368,g13385,g13390,g13395,g13477,g13479,g13480,g13481,g13483,g13484,
    g13485,g13486,g13487,g13488,g13489,g13490,g13491,g13492,g13493,g13496,
    g13498,g13499,g13500,g13502,g13503,g13504,g13505,g13506,g13513,g13515,
    g13516,g13517,g13527,g13609,g13619,g13623,g13625,g13631,g13634,g13636,
    g13642,g13643,g13645,g13646,g13648,g13654,g13655,g13656,g13671,g13672,
    g13674,g13675,g13676,g13701,g13702,g13703,g13704,g13705,g13738,g13739,
    g13740,g13755,g13787,g13788,g13789,g13790,g13796,g13815,g13816,g13818,
    g13824,g13833,g13834,g13835,g13837,g13839,g13845,g13846,g13847,g13851,
    g13853,g13854,g13855,g13860,g13862,g13870,g13871,g13878,g13880,g13884,
    g13892,g13900,g13902,g13904,g13905,g13913,g13914,g13933,g13941,g13943,
    g13944,g13952,g13953,g13969,g13970,g13989,g13997,g13998,g14006,g14007,
    g14022,g14023,g14039,g14040,g14059,g14067,g14097,g14098,g14113,g14114,
    g14130,g14131,g14143,g14182,g14212,g14213,g14228,g14229,g14297,g14327,
    g14328,g14336,g14419,g14690,g14724,g14752,g14767,g13245,g14773,g14884,
    g14894,g14956,g14957,g14958,g14975,g15020,g15030,g15031,g15046,g15047,
    g15064,g15093,g15094,g15104,g15105,g15126,g15127,g15142,g15143,g15160,
    g15171,g15172,g15173,g15178,g15196,g15197,g15218,g15219,g15234,g15235,
    g15243,g15244,g15245,g15246,g15247,g15257,g15258,g15259,g15264,g15282,
    g15283,g15304,g15305,g15320,g15321,g15324,g15325,g15335,g15336,g15337,
    g15338,g15339,g15349,g15350,g15351,g15356,g15374,g15375,g15388,g15389,
    g15391,g15392,g15402,g15403,g15407,g15410,g15411,g15421,g15422,g15423,
    g15424,g15425,g15435,g15436,g15437,g15442,g15452,g15453,g15459,g15460,
    g15470,g15475,g15476,g15486,g15487,g15491,g15494,g15495,g15505,g15506,
    g15507,g15508,g15509,g15519,g15520,g15526,g15527,g15545,g15546,g15556,
    g15561,g15562,g15572,g15573,g15577,g15580,g15581,g15591,g15592,g15593,
    g15594,g15595,g15604,g15605,g15623,g15624,g15634,g15639,g15640,g15650,
    g15651,g15658,g15666,g15670,g15671,g15680,g15681,g15699,g15700,g15710,
    g15717,g15725,g15729,g15730,g15739,g15740,g15753,g15754,g15755,g15765,
    g15769,g15770,II22028,g15780,g15781,g15793,g15801,g15802,g15817,g15828,
    g15829,g15840,g15852,II22136,g15902,g15998,g16003,g16004,g16008,g16009,
    g16010,g16015,g16016,g16017,g16018,g16019,g16028,g16029,g16030,g16031,
    g16032,g16033,g16045,g16046,g16047,g16048,g16049,g16050,g16051,g16052,
    g16066,g16067,g16068,g16069,g16070,g16071,g16072,g16073,g16074,g16089,
    g16100,g16101,g16102,g16103,g16104,g16105,g16106,g16107,g16108,g16111,
    g16112,g16119,g16127,g16133,g16134,g16135,g16136,g16137,g16138,g16139,
    g16140,g16141,g16153,g16158,g16159,g16160,g16161,g16162,g16163,g16170,
    g16178,g16182,g16183,g16184,g16185,g16186,g16187,g16188,g16198,g16199,
    g16200,g16211,g16212,g16217,g16218,g16219,g16220,g16221,g16222,g16229,
    g16237,g16238,g16239,g16240,g16241,g16242,g16251,g16252,g16253,g16262,
    g16263,g16264,g16265,g16276,g16277,g16282,g16283,g16284,g16285,g16286,
    g16288,g16289,g16290,g16291,g16298,g16299,g16300,g16301,g16309,g16310,
    g16311,g16312,g16321,g16322,g16323,g16324,g16335,g16336,g16342,g16343,
    g16344,g16345,g16347,g16348,g16349,g16350,g16356,g16357,g16358,g16359,
    g16367,g16368,g16369,g16370,g16379,g16380,g16381,g16382,g16383,g16385,
    g16386,g16387,g16388,g16389,g16390,g16391,g16392,g16393,g16394,g16400,
    g16401,g16402,g16403,g16411,g16413,g16414,g16415,g16416,g16417,g16418,
    g16419,g16420,g16421,g16422,g16423,g16424,g16425,g16426,g16427,g16428,
    g16429,g16430,g16431,g16432,g16438,g16443,g16444,g16445,g16447,g16448,
    g16449,g16450,g16451,g16452,g16453,g16454,g16455,g16456,g16457,g16458,
    g16459,g16460,g16461,g16462,g16505,g16513,g16527,g16535,g16558,g16590,
    g16607,g16625,g16639,g16650,g16850,g16855,g16856,g16859,g16864,g16865,
    g16879,g16894,g16907,g16908,g16909,g16923,g16938,g16939,g16953,g16964,
    g16966,g16967,g16968,g16969,g16970,g16984,g16987,g16988,g16989,g16990,
    g16991,g16993,g16994,g16997,g16998,g16999,g17001,g17015,g17017,g17018,
    g17021,g17022,g17023,g17028,g17031,g17045,g17047,g17048,g17055,g17056,
    g17062,g17065,g17079,g17081,g17082,g17084,g17090,g17091,g17097,g17100,
    g17114,g17116,g17117,g17122,g17128,g17129,g17135,g17138,g17143,g17144,
    g17149,g17155,g17156,g17161,g17166,g17167,g17172,g17176,g17181,g17182,
    g17193,g17268,g17301,g17339,g17352,g17353,g17381,g17382,g17393,g17395,
    g17396,g17397,g17398,g17408,g17409,g17428,g17446,g17447,g17448,g17449,
    g17450,g17460,g17461,g17462,g17463,g17464,g17474,g17475,g17485,g17486,
    g17506,g17508,g17509,g17510,g17526,g17527,g17528,g17529,g17530,g17540,
    g17541,g17542,g17543,g17544,g17554,g17555,g17556,g17576,g17577,g17578,
    g17597,g17598,g17599,g17600,g17616,g17617,g17618,g17619,g17620,g17630,
    g17631,g17632,g17633,g17634,g17635,g17636,g17652,g17653,g17654,g17673,
    g17674,g17675,g17694,g17695,g17696,g17697,g17713,g17714,g17715,g17716,
    g17717,g17718,g17719,g17734,g17735,g17736,g17737,g17752,g17753,g17754,
    g17773,g17774,g17775,g17794,g17795,g17796,g17797,g17798,g17812,g17813,
    g17814,g17824,g17835,g17836,g17837,g17838,g17853,g17854,g17855,g17874,
    g17875,g17876,g17877,g17900,g17901,g17902,g17912,g17924,g17925,g17926,
    g17936,g17947,g17948,g17949,g17950,g17965,g17966,g17967,g17989,g17990,
    g18011,g18012,g18013,g18023,g18035,g18036,g18037,g18047,g18058,g18059,
    g18060,g18061,g18062,g18088,g18106,g18107,g18128,g18129,g18130,g18140,
    g18152,g18153,g18154,g18164,g18165,g18169,g18204,g18222,g18223,g18244,
    g18245,g18246,g18256,g18311,g18329,g18330,g18333,g18404,II24619,g18547,
    II24689,g18597,II24738,g18629,II24758,g18638,g18645,g18647,g18648,g18649,
    g18650,g18651,g18652,g18653,g18654,g18655,g18665,g18666,g18667,g18668,
    g18688,g18689,g18690,g18717,g18718,g18753,g18982,g18990,g18994,g18997,
    g19007,g19010,g19063,g19079,g19080,g19087,g17215,g19088,g19089,g19090,
    g19092,g19093,g17218,g19094,g19095,II25280,g19097,g19099,g19100,g17220,
    g19101,g19102,II25291,g19104,g19106,g19107,g17223,g19108,II25300,g19109,
    g19111,g19112,II25311,g19116,g19117,g19124,g19131,g19142,g17159,g19143,
    g17174,g19146,g17191,g19148,g17202,g19150,g19155,g19161,g19166,g19228,
    g16662,g19236,g16935,g19241,g19248,g19252,g19254,g19260,g19267,g19282,
    g19284,g19285,g19289,g19303,g19307,g19316,g19317,g19320,g19324,g19328,
    g19347,g19351,g19355,g19356,g19381,g19385,g19413,g19449,g19476,g19499,
    g19520,g19531,g19540,g19541,g19544,g19545,g19547,g19548,g19549,g19551,
    g19552,g16829,g19553,g19554,g19555,g19557,g19558,g19559,g19560,g19561,
    g19562,g19564,g19565,g19566,g19567,g19568,g19569,g19570,g19571,g19572,
    g19574,g19575,g19576,g19584,g19585,g19586,g19587,g19588,g19589,g19590,
    g19591,g19592,g19593,g19594,g19597,g19598,g19599,g19600,g19601,g19602,
    g19603,g19604,g19605,g19606,g19614,g19615,g19616,g19617,g19618,g19619,
    g19620,g19621,g19623,g19624,g19625,g19626,g19627,g19628,g19629,g19630,
    g19631,g19632,g19633,g19634,g19635,g19636,g19637,g19638,g19639,g19647,
    g19648,g19649,g19650,g19651,g19653,g19654,g19655,g19656,g19660,g19661,
    g19662,g19663,g19664,g19665,g19666,g19667,g19668,g19669,g19670,g19671,
    g19672,g19673,g19674,g19675,g19676,g19677,g19678,g19679,g19687,g19688,
    g19691,g16841,g19692,g19693,g19694,g19695,g19697,g19698,g19699,g19700,
    g19701,g19702,g19703,g19704,g19708,g19709,g19710,g19711,g19712,g19713,
    g19714,g19715,g19716,g19717,g19718,g19719,g19720,g19721,g19722,g19723,
    g19724,g19726,g16847,g19727,g19728,g19729,g19730,g19731,g19732,g19733,
    g19734,g19735,g19736,g19737,g19738,g19739,g19741,g19742,g19743,g19744,
    g19745,g19746,g19747,g19748,g19752,g19753,g19754,g19755,g19756,g19757,
    g19758,g19759,g19760,g19761,g19764,g19765,g19766,g19767,g19768,g19769,
    g19770,g19771,g19772,g19773,g19774,g19775,g19776,g19777,g19778,g19779,
    g19780,g19781,g19782,g19784,g19785,g19786,g19787,g19788,g19789,g19790,
    g19791,g19795,g19796,g19797,II26240,g19799,g19802,g19803,g19804,g19805,
    g19806,g19807,g19808,g19809,g19810,g19811,g19812,g19813,g19814,g19815,
    g19816,g19817,g19818,g19819,g19820,g19821,g19822,g19823,g19824,g19826,
    g19827,g19828,g19829,g19836,g19837,g19839,g19840,g19841,II26282,g19842,
    II26285,g19843,g19846,g19847,g19848,g19849,g19850,g19851,g19852,g19853,
    g19854,g19855,g19856,g19857,g19858,g19859,g19860,g19861,g19862,g19863,
    g19864,g19868,g16498,g19869,g19870,II26311,g19871,g19872,g19873,g19874,
    II26317,g19875,II26320,g19876,g19879,g19880,g19881,g19882,g19883,g19884,
    g19885,g19886,g19887,g19888,g19889,g19895,g19899,g16520,g19900,g19901,
    II26348,g19902,g19903,g19904,g19905,II26354,g19906,II26357,g19907,g19910,
    g19911,g19912,g19913,g19914,g19920,g19924,g16551,g19925,g19926,II26377,
    g19927,g19928,g19929,g19930,II26383,g19931,g19932,g19935,g19939,g16583,
    g19940,g19941,II26396,g19942,g19943,g19944,g19949,g19952,g19953,II26416,
    g18553,g18491,g18431,g19970,g18354,g18276,g19971,g19976,II26432,g18277,
    g18189,g18090,g19982,g17992,g17913,g19983,II26440,g18603,g18555,g18504,
    g20000,g18449,g18369,g20001,g20006,g20011,g20012,g20013,g20014,II26464,
    g18370,g18296,g18206,g20020,g18109,g18024,g20021,II26472,g18635,g18605,
    g18568,g20038,g18522,g18464,g20039,g20044,g20048,g20049,g20050,g20051,
    g20052,g20053,II26500,g18465,g18389,g18313,g20062,g18225,g18141,g20063,
    II26508,g18644,g18637,g18618,g20080,g18586,g18537,g20081,g20084,g20085,
    g20086,g20087,g20088,g20089,g20090,g20091,g20092,II26525,g20093,II26528,
    g20094,II26541,g18538,g18484,g18406,g20103,g18332,g18257,g20104,g20106,
    g20107,g20108,g20109,g20110,g20111,g20112,g20113,g20114,g20115,II26558,
    g20116,II26561,g20117,II26564,g20118,II26567,g20119,g20131,g20132,g20133,
    g20134,g20135,g20136,g20137,g20138,g20139,g20144,g16679,g20145,II26590,
    g20146,II26593,g20147,II26596,g20148,II26599,g20149,g20156,g20157,g20158,
    g20159,g20160,g20161,g20162,II26615,g20177,g20182,g16705,g20183,II26621,
    g20184,II26624,g20185,II26627,g20186,II26630,g20187,g20188,g20189,g20190,
    g20191,g20192,II26639,g20197,II26645,g20211,g20216,g16736,g20217,II26651,
    g20218,II26654,g20219,g20220,g20221,g20222,II26661,g20227,II26667,g20241,
    g20246,g16778,g20247,g20248,g20249,II26676,g20254,II26682,g20268,g20270,
    g20271,g20272,II26690,g20277,II26695,g20280,g20282,g20283,g20284,g20285,
    II26708,g20291,g20293,g20294,II26726,g20307,g20309,II26745,g20326,g20460,
    g20472,g20480,g20486,g20492,g20499,g20502,g20503,g17507,g20506,g20512,
    g20525,g20538,g20640,g20647,g20665,g20809,g20826,g20836,g20840,g21049,
    g21067,g21068,g21077,g21078,g21085,g21086,g21091,g21092,g21097,g21098,
    g21103,g21107,g21111,g21112,g21121,g20054,g21122,g21123,g21124,g21128,
    g21129,II27695,g19318,g19300,g19286,g21136,g19271,g19261,g21137,g21138,
    g21140,g20095,g21141,g21142,g21143,II27711,g19262,g19414,g19386,g21152,
    g19357,g19334,g21153,g21154,g21155,II27717,g19345,g19321,g19304,g21156,
    g19290,g19276,g21157,g21158,g21160,g20120,g21161,g21162,g21163,II27733,
    g19277,g19451,g19416,g21172,g19389,g19368,g21173,g21174,g21175,II27739,
    g19379,g19348,g19325,g21176,g19308,g19295,g21177,g21178,g21180,g20150,
    g21181,g21182,g21188,II27755,g19296,g19478,g19453,g21192,g19419,g19400,
    g21193,g21194,g21195,II27761,g19411,g19382,g19352,g21196,g19329,g19313,
    g21197,g21198,g21203,II27772,g19314,g19501,g19480,g21207,g19456,g19430,
    g21208,g21209,g21210,g21218,g21226,g21229,g21234,g21243,g21245,g20299,
    g21251,g21252,g21254,g20318,g21259,g21260,g21262,g20337,g21267,g21268,
    g21270,g20357,g21276,g21277,g21283,g21284,g21290,g21291,g21292,g21298,
    g21299,g21300,g21301,g21302,g21303,g21304,g21305,g21306,g21307,g21308,
    g21309,g21310,g21311,g21312,g21313,g21314,g21315,g21319,g21320,g21321,
    g21322,g21323,g21324,g21325,g21326,g21328,g21329,g21330,g21334,g21335,
    g21336,g21337,g21338,g21339,g21340,g21341,g21342,g21343,g21344,g21345,
    g21349,g21350,g21351,g21352,g21353,g21354,g21355,g21356,g21357,g21360,
    g21361,g21362,g21363,g21367,g21368,g21369,g21370,g21371,g21372,g21373,
    g21374,g21375,g21378,g21379,g21380,g21381,g21388,g21389,g21390,g21391,
    g21392,g21393,g21394,g21395,g21396,g21397,g21398,g21401,g21402,g21403,
    g21410,g21411,g21412,g21413,g21414,g21418,g21419,g21420,g21421,g21422,
    g21423,g21424,g21425,g21428,g21438,g21439,g21440,g21444,g21445,g21446,
    g21447,g21448,g21452,g21453,g21454,g21455,g21456,g21476,g21480,g21481,
    g21482,g21486,g21487,g21488,g21489,g21490,g21494,g21497,g21517,g21521,
    g21522,g21523,g21527,II28068,g21553,II28096,g21564,II28103,g21589,g21593,
    II28126,g21597,II28133,g21610,g21611,g21622,II28155,g21626,II28162,g21635,
    g21639,g21650,II28181,g21654,g21658,g21666,g21670,g21681,g21687,g21695,
    g21699,g21707,g21723,g21731,g21735,g21749,g21757,g21758,g21773,g21805,
    g21812,g21818,g21822,g21891,g21892,g19288,g21899,g21900,g19306,g21906,
    g21911,g21912,g19327,g21913,g21920,g21925,g21926,g19354,g21931,g21938,
    g21990,g22004,g22015,g22020,II28582,g19141,g21133,g21116,g21104,g21095,
    g21084,II28594,g21167,g21147,g21134,g21117,g21105,g21096,II28609,g21183,
    g21168,g21148,g21135,g21118,g21106,g22187,g22196,g22201,g22202,g22206,
    g22207,g22208,g22211,g22214,g22215,g22220,g22223,g22224,g22228,g22229,
    g22235,g22238,g22244,g22245,g22250,g22254,g22255,g22264,g22265,g22270,
    g22272,g22273,g22281,g22282,g22285,g22289,g22291,g22292,g22305,g22309,
    g22311,g22312,g22333,g22337,g22340,g22358,g22363,g22383,g22398,g22483,
    g22515,g22516,g22517,g22526,g22546,g22555,g22556,g22557,g22566,g22577,
    g22581,g22587,g22595,g22596,g22597,g22606,g22607,g22610,g22614,g22618,
    g22624,g22632,g22633,g22634,g22637,g20841,g22638,g22643,g22646,g22650,
    g22654,g22660,g22665,g20920,g22666,g22667,g22674,g22679,g22682,g22686,
    g22690,g22699,g22700,g22701,g22707,g22714,g22719,g22722,g22726,g22727,
    g22732,g22738,g22745,g22754,g22759,g22764,g22770,g22788,g22793,g22798,
    g22804,g22830,g22835,g22841,g22842,g22869,g22874,g22906,g22984,g23104,
    g23106,g23118,g23119,g23127,g23128,g23138,g23139,g23409,g23414,g23419,
    g22755,g23423,g23428,g22789,g23432,g23434,g22831,g23440,g22870,g23451,
    g23458,g23462,g23467,g23471,g23476,g23483,g23484,g23494,g23496,g23510,
    g23512,g23525,g23527,g23536,g23538,g23544,g23547,g23550,g23551,g23552,
    g23554,g23558,g23559,g23560,g23563,g23564,g23565,g23567,g23571,g23572,
    g23573,g23577,g23578,g23579,g23582,g23583,g23584,g23586,g23590,g23591,
    g23592,g23593,g22845,g23598,g23599,g23600,g23604,g23605,g23606,g23609,
    g23610,g23611,g23615,g23616,g23617,g22810,g23618,g22608,g23622,g23623,
    g23624,g23625,g22880,g23630,g23631,g23632,g23636,g23637,g23638,g23639,
    g23643,g23659,g22784,g23664,g23665,g23666,g22851,g23667,g22644,g23671,
    g23672,g23673,g23674,g22915,g23679,g23680,g23681,g23686,g23687,g22668,
    g23689,g23693,g23709,g22826,g23714,g23715,g23716,g22886,g23717,g22680,
    g23721,g23722,g23723,g23724,g22940,g23726,g23734,g23735,g23740,g23741,
    g22708,g23743,g23747,g23763,g22865,g23768,g23769,g23770,g22921,g23771,
    g22720,g23772,g23776,g23777,g23778,g23789,g23790,g23795,g23796,g22739,
    g23798,g23802,g23818,g22900,g23820,g23822,g23824,g23825,g23829,g23830,
    g23831,g23842,g23843,g23848,g23849,g22771,g23851,g23852,g19179,g23854,
    g23855,g23857,g23859,g23860,g23864,g23865,g23866,g23877,g23878,g23886,
    g23888,g23889,g23891,g23893,g23894,g23898,g23899,g23900,g23904,g23907,
    g23909,g23910,g23912,g23914,g23915,g23917,g23939,g23941,g23942,g23944,
    g23971,g23972,g24029,g24211,g24217,g24221,g24224,g24229,g24236,g24241,
    g24246,g24247,g24253,g24256,g24427,g24429,g24431,g24432,g24433,g24435,
    g24436,g24437,g24439,g24440,g24441,g23545,g21119,g21227,g24529,g24540,
    g24541,g24542,g24550,g24552,g24553,g24554,g24559,g24561,g24563,g24564,
    g24565,g24569,g24571,g24573,g24574,g24578,g24580,g24585,g24590,g24591,
    g24595,g24596,g24603,g24604,g24610,g24611,g24644,g24664,g24683,g24700,
    g24745,g15454,g24746,g24747,g24748,g24749,g15540,g24750,g24751,g24752,
    g24754,g24755,g24757,g24758,g15618,g24759,g24760,g24761,g24762,g24767,
    g24768,g24769,g24772,g24773,g24774,g24775,g15694,g24776,g24777,g24779,
    g24780,g24781,g24788,g24789,g24790,g24792,g24793,g24794,g24795,g24232,
    g24796,g24798,g24799,g24802,g24803,g24804,g24809,g24810,g24811,g24813,
    g24818,g24821,g24822,g24824,g24825,g24826,g24831,g24100,g24838,g24840,
    g24841,g24843,g24846,g24109,g24853,g24855,g24858,g24861,g24126,g24867,
    g24869,g24870,g24874,g24876,g24145,g24878,g24881,g24882,g24884,g24885,
    g24888,g24898,g24899,g24901,g24902,g24905,g24906,g24907,g24908,g24921,
    g24922,g24924,g24938,g24964,g24974,g25086,g25102,g25117,g25128,g25178,
    g24623,g25181,g24636,g25182,g24681,g25184,g24694,g25187,g24633,g25188,
    g24652,g25192,g24711,g25193,g24653,g25196,g24672,g25198,g24691,g25269,
    g25277,g25278,g25281,g25282,g25286,g25287,g25289,g25290,g25294,g25295,
    g25299,g25300,g25304,g25309,g25310,g25318,g24682,g25321,g25075,g25328,
    g25334,g25337,g25342,g25346,g25348,g25351,g25356,g25360,g25362,g25365,
    g25371,g25375,g25377,g25388,g25392,g25453,g25457,g25461,g25466,g25470,
    g24479,g25475,g25482,g24480,g25483,g24481,g25487,g24485,g25505,g25506,
    g25513,g24487,g25514,g24488,g25518,g24489,g25552,g25553,g25560,g24494,
    g25561,g24495,g25565,g24496,g25618,g25619,g25626,g24504,g25627,g24505,
    g25628,g21008,g25629,g25697,g25881,g25951,g24800,g25953,g24783,g25957,
    g24782,g25961,g24770,g25963,g24756,g25968,g24871,g25972,g24859,g25973,
    g24847,g25975,g24606,g25977,g24845,g25978,g24836,g25980,g24663,g25981,
    g24819,g26023,g26024,g26026,g26027,g25418,g26028,g26029,g26030,g25429,
    g26032,g26033,g26034,g26035,g25523,g26036,g26038,g25589,g26039,g25668,
    g26040,g25745,g26051,g26052,g25941,g26053,g26054,g25944,g26060,g25943,
    g26061,g26062,g25947,g26067,g25946,g26068,g26069,g25949,g26074,g25948,
    g26075,g26080,g25950,g26082,g26085,g26091,g26157,g26158,g26163,g26166,
    g26171,g26186,g26188,g26207,g26212,g26213,g26231,g26233,g26234,g26235,
    g26236,g26243,g26244,g26257,g26258,g26259,g26260,g25254,g26261,g26262,
    g26263,g26268,g26269,g26270,g26271,g26278,g26279,g26288,g26289,g26290,
    g26291,g26292,g26293,g26298,g26299,g26300,g26301,g25258,g26302,g26303,
    g26307,g26309,g26310,g26311,g26312,g26316,g26317,g26318,g26319,g26324,
    g26325,g26326,g26332,g26333,g26334,g26335,g26339,g26340,g26342,g26343,
    g26344,g26345,g25261,g26346,g26347,g26348,g26350,g26351,g26352,g26353,
    g26357,g26361,g26362,g26363,g26365,g26366,g26371,g26372,g26373,g26379,
    g26380,g26381,g26382,g26383,g26384,g26386,g26387,g26388,g26389,g25264,
    g26390,g26391,g26392,g26396,g26397,g26400,g26404,g26405,g26406,g26408,
    g26409,g26414,g26415,g26416,g26422,g26423,g26424,g26425,g26426,g26427,
    g26432,g26437,g26438,g26441,g26445,g26446,g26447,g26449,g26450,g26455,
    g26456,g26457,g26464,g26469,g26470,g26473,g26477,g26478,g26479,g26488,
    g26493,g26494,g26504,g26663,g26668,g26673,g12431,g26674,g26754,g26755,
    g26083,g26756,g26113,g26758,g16614,g26759,g26356,g26760,g26137,g26761,
    g26154,g26763,g26764,g16632,g26765,g26399,g26766,g26767,g26087,g26768,
    g26440,g26769,g26770,g26059,g26771,g26773,g26145,g26774,g26472,g26775,
    g26099,g26777,g26066,g26778,g26780,g26119,g26783,g26073,g26784,g26787,
    g26129,g26790,g26079,g26791,g26794,g26143,g26797,g26148,g26829,g26833,
    g26842,g26845,g26851,g26853,g26860,g26866,g26955,g26958,g26961,g26962,
    g26963,g26965,g23320,g26966,g26967,g26968,g26969,g26970,g21976,g26971,
    g23325,g26972,g26973,g26977,g26978,g26979,g23331,g26980,g23360,g26981,
    g26982,g21983,g26984,g23335,g26985,g26986,g26993,g26994,g26995,g21991,
    g26996,g26997,g22050,g26998,g26999,g27000,g23340,g27001,g23364,g27002,
    g27003,g21996,g27004,g23344,g27005,g27006,g27007,g27008,g27009,g23368,
    g27016,g27017,g27018,g22005,g27019,g27020,g22069,g27021,g27022,g27023,
    g23349,g27024,g23372,g27025,g27026,g22009,g27027,g27028,g27029,g27030,
    g22083,g27031,g27032,g27033,g27034,g27035,g23377,g27042,g27043,g27044,
    g22016,g27045,g27046,g22093,g27047,g27048,g27049,g23353,g27050,g23381,
    g27052,g27053,g27054,g27055,g27056,g27057,g27058,g22108,g27059,g27060,
    g27061,g27062,g27063,g23388,g27070,g27071,g27072,g22021,g27073,g27074,
    g22118,g27076,g27077,g27079,g27080,g27081,g27082,g27083,g27084,g27085,
    g22134,g27086,g27087,g27088,g27089,g27090,g23395,g27091,g27092,g27093,
    g27095,g27096,g27097,g27098,g27099,g27100,g27101,g22157,g27103,g27104,
    g27105,g27107,g27108,g27109,g27110,g27111,g27112,g27115,g27178,g26110,
    g27181,g16570,g27182,g26151,g27185,g26126,g27187,g16594,g27240,g26905,
    g27241,g26934,g27242,g27244,g26914,g27245,g26877,g27246,g26988,g27247,
    g27011,g27248,g27037,g27249,g27065,g27355,g27356,g27358,g27359,g27364,
    g27365,g27370,g27371,g27372,g27394,g27396,g27407,g27409,g27425,g27427,
    g27446,g27448,g27495,g23945,g27509,g27516,g23974,g27530,g27534,g27541,
    g24004,g27552,g27554,g27561,g24038,g27568,g27570,g27578,g27656,g27657,
    g27659,g27660,g27661,g27666,g27671,g26885,g27673,g27679,g27680,g27681,
    g27719,g27496,g27720,g27481,g27721,g27579,g27723,g27464,g27725,g27532,
    g27726,g27531,g27727,g27414,g27728,g27564,g27729,g27435,g27730,g27454,
    g27731,g27470,g27732,g27492,g27733,g27513,g27734,g27538,g27737,g27558,
    g27770,g27772,g27773,g27774,g27775,g27779,g27783,g27790,g27904,g27908,
    g27909,g27913,g27914,g27915,g27922,g27923,g27924,g27926,g27931,g27935,
    g27936,g27938,g27945,g27949,g27951,g27963,g27968,g27970,g27984,g27985,
    g27991,g28008,g28009,g28015,g28027,g28028,g28035,g28036,g28042,g28050,
    g28051,g28057,g28058,g28065,g28066,g28073,g28079,g28080,g28086,g28087,
    g28094,g28098,g28104,g28105,g28111,g28112,g28116,g28122,g28123,g28127,
    g28171,g28176,g28188,g28193,g27573,g28319,g27855,g28320,g27854,g28322,
    g27937,g28323,g27838,g28324,g27810,g28326,g27865,g28327,g27900,g28329,
    g27823,g28330,g27864,g28331,g27802,g28332,g27883,g28333,g27882,g28334,
    g27842,g28335,g27814,g28336,g27896,g28337,g28002,g28338,g28029,g28339,
    g28059,g28340,g28088,g28373,g28376,g28378,g28379,g27868,g28380,g28381,
    g28157,g28383,g28385,g28387,g28389,g28396,g28398,g28399,g28401,g28402,
    g28404,g28405,g28407,g28408,g28411,g28412,g28416,g28422,g28423,g28424,
    g28426,g28427,g28428,g28429,g28430,g28431,g28433,g28434,g28435,g28436,
    g28438,g28439,g28440,g28441,g28442,g28444,g28445,g28446,g28448,g28450,
    g28451,g28452,g28453,g28454,g28456,g28457,g28459,g28460,g28462,g28463,
    g28464,g28465,g28466,g28468,g28469,g28471,g28472,g28474,g28475,g28476,
    g28477,g28478,g28479,g28480,g28481,g28484,g28485,g28486,g28487,g28492,
    g28493,g28494,g28497,g28657,g27925,g28659,g27917,g28660,g27916,g28662,
    g27911,g28663,g27906,g28664,g27997,g28665,g27827,g28666,g27980,g28667,
    g27964,g28669,g27897,g28670,g27798,g28671,g27962,g28672,g27950,g28707,
    g12436,g28708,g28392,g28709,g28400,g28710,g28403,g28711,g28415,g28712,
    g28406,g28713,g28410,g28714,g28394,g28715,g28414,g28716,g28449,g28717,
    g28461,g28718,g28473,g28719,g28482,g28722,g28523,g28724,g28551,g28726,
    g28578,g28729,g28606,g28834,g28836,g28838,g28840,g28841,g27834,g28843,
    g28844,g27850,g28846,g28847,g28848,g27875,g28849,g28850,g28851,g27892,
    g28852,g28853,g28854,g28880,g28881,g28892,g28893,g28897,g28898,g28909,
    g28910,g28914,g28915,g28919,g28923,g28931,g28935,g28936,g28940,g28944,
    g28948,g28949,g28958,g28962,g28966,g28970,g28971,g28986,g28996,g28997,
    g29022,g29130,g28397,g29174,g29031,g29175,g29009,g29176,g29097,g29180,
    g28982,g29183,g29064,g29186,g29063,g29188,g29083,g29196,g29200,g29203,
    g29208,g29211,g29217,g29220,g29225,g29229,g29232,g29233,g29234,g29235,
    g29236,g29238,g29239,g29240,g29241,g29242,g29243,g29248,g29251,g29252,
    g29255,g29256,g29257,g29259,g29260,g29261,g29262,g29263,g29264,g29284,
    g29001,g29289,g29030,g29294,g29053,g29300,g29072,g29302,g29026,g29310,
    g28978,g29312,g29049,g29320,g29088,g29321,g29008,g29323,g29068,g29329,
    g29096,g29330,g29038,g29332,g29080,g29336,g29045,g29337,g29103,g29338,
    g29060,g29341,g29062,g29342,g29107,g29344,g29076,g29346,g29087,g29411,
    g29090,g29464,g29465,g29466,g29265,g29467,g29340,g29468,g29343,g29469,
    g29345,g29470,g29347,g29471,g29472,g29473,g29474,g29475,g29476,g29477,
    g29478,g29479,g29480,g29481,g29482,g29483,g29484,g29485,g29486,g29487,
    g29488,g29489,g29490,g29502,g29518,g28728,g29520,g28731,g29521,g28733,
    g29522,g27735,g29523,g28737,g29524,g28739,g29525,g29195,g29526,g27741,
    g29527,g28748,g29528,g28750,g29529,g29199,g29531,g29202,g29532,g27746,
    g29533,g28762,g29534,g29206,g29536,g29207,g29538,g29210,g29539,g27754,
    g29540,g26041,g29541,g29214,g29543,g29215,g29545,g29216,g29547,g29219,
    g29548,g28784,g29549,g26043,g29550,g29222,g29553,g29223,g29555,g29224,
    g29557,g28789,g29558,g28790,g29559,g26045,g29560,g29227,g29562,g29228,
    g29564,g28794,g29565,g28795,g29566,g26047,g29567,g29231,g29572,g28802,
    g29573,g28803,g29575,g28813,g29607,g29610,g29614,g29615,g29619,g29622,
    g29624,g29625,g29626,g29790,g29792,g29793,g29810,g29748,g29811,g29703,
    g29812,g29762,g29813,g29760,g29814,g29728,g29815,g29727,g29816,g29759,
    g29817,g29709,g29818,g29732,g29819,g29751,g29820,g29717,g29821,g29731,
    g29822,g29705,g29827,g29741,g29828,g29740,g29833,g29725,g29834,g29713,
    g29839,g29747,g29909,g29735,g29910,g29779,g29942,g29771,g29944,g29782,
    g29945,g29773,g29946,g29778,g29947,g29785,g29948,g29775,g29949,g29781,
    g29950,g29788,g29951,g29777,g29952,g29784,g29953,g29791,g29954,g29770,
    g29955,g29787,g29956,g29780,g29957,g29772,g29958,g29783,g29959,g29774,
    g29960,g29786,g29961,g29776,g29962,g29789,g29963,g29758,g29964,g29757,
    g29965,g29756,g29966,g29755,g29967,g29754,g29968,g29765,g29969,g29721,
    g29970,g29764,g29971,g29763,g29980,g29981,g29982,g29983,g29984,g29985,
    g29986,g29987,g29988,g29989,g29990,g29991,g29992,g12441,g29993,g29994,
    g29995,g29996,g29997,g29918,g29998,g29922,g29999,g29924,g30000,g29930,
    g30001,g30002,g30003,g30004,g29926,g30005,g30006,g29928,g30007,g30008,
    g29919,g30009,g29929,g30077,g30079,g30080,g30081,g30082,g30083,g30085,
    g30086,g30087,g30088,g30089,g30090,g30091,g30092,g30093,g30094,g30095,
    g30096,g30097,g30098,g30099,g30100,g30101,g30102,g30103,g30104,g30105,
    g30106,g30107,g30108,g30109,g30110,g30111,g30112,g30113,g30114,g30115,
    g30116,g29921,g30117,g30118,g30123,g30070,g30127,g30065,g30128,g30062,
    g30129,g30071,g30131,g30059,g30132,g30068,g30133,g30067,g30138,g30069,
    g30216,g30217,g30218,g30219,g30220,g30221,g30222,g30223,g30224,g30225,
    g30226,g30227,g30327,g30330,g30333,g30334,g30337,g30340,g30345,g30348,
    g30351,g30352,g30355,g30361,g30364,g30367,g30372,g30228,g30374,g30387,
    g30388,g30389,g30390,g30391,g30392,g30393,g30394,g30395,g30396,g30397,
    g30398,g30407,g30409,g30410,g30411,g30436,g30437,g30438,g30440,g30441,
    g30442,g30444,g30445,g30447,g30448,g30449,g30451,g30452,g30453,g30454,
    g30457,g30458,g30460,g30461,g30462,g30464,g30465,g30467,g30469,g30472,
    g30473,g30475,g30476,g30477,g30478,g30481,g30484,g30486,g30489,g30490,
    g30492,g30495,g30496,g30499,g30502,g30504,g30696,g30697,g30698,g30728,
    g30605,g30735,g30629,g30736,g30584,g30743,g30610,g30744,g30609,g30750,
    g30593,g30754,g30614,g30755,g30632,g30757,g30601,g30758,g30613,g30759,
    g30588,g30760,g30622,g30761,g30621,g30762,g30608,g30763,g30597,g30764,
    g30628,g30766,g30617,g30916,g30785,g30917,g12446,g30918,g30780,g30919,
    g30786,g30920,g30787,g30921,g30791,g30922,g30788,g30923,g30789,g30924,
    g30783,g30925,g30790,g30944,g30935,g30945,g30931,g30946,g30930,g30947,
    g30936,g30948,g30929,g30949,g30933,g30950,g30932,g30951,g30934,g30953,
    g30952,g9144,g10778,g12377,g12407,g12886,g12926,g12955,g12984,g16539,
    g16571,g16595,g16615,g19181,g17729,g17979,g19186,g18419,g17887,g19187,
    g19188,g17830,g18096,g19191,g17807,g19192,g18183,g18270,g19193,g18492,
    g17998,g19194,g19195,g17942,g18212,g19200,g18346,g18424,g19201,g19202,
    g17919,g19203,g18290,g18363,g19204,g18556,g18115,g19205,g19206,g18053,
    g18319,g19209,g18079,g19210,g19211,g18441,g18497,g19212,g19213,g18030,
    g19214,g18383,g18458,g19215,g18606,g18231,g19216,g19221,g19222,g18195,
    g19223,g19224,g18514,g18561,g19225,g19226,g18147,g19227,g18478,g18531,
    II25477,g17024,g17000,g16992,g19230,g16985,g16965,g19231,g19232,g18302,
    g19233,g19234,g18578,g18611,g19235,II25495,g17158,g17137,g17115,g19240,
    g17083,g17050,g19242,II25500,g17058,g17030,g17016,g19243,g16995,g16986,
    g19244,g19245,g18395,g19246,g19250,II25516,g17173,g17160,g17142,g19253,
    g17121,g17085,g19255,II25521,g17093,g17064,g17046,g19256,g17019,g16996,
    g19257,g19263,g19264,II25549,g17190,g17175,g17165,g19266,g17148,g17123,
    g19268,II25554,g17131,g17099,g17080,g19269,g17049,g17020,g19275,g19278,
    g19279,II25588,g17201,g17192,g17180,g19281,g17171,g17150,g19283,g19294,
    g19297,g19298,g19312,g19315,g19333,g19450,g19477,g19500,g19503,g19521,
    g19522,g19532,g19542,II26429,g19981,II26455,g20015,II26461,g20019,II26491,
    g20057,II26497,g20061,II26532,g20098,II26538,g20102,II26571,g20123,g21120,
    g21139,g21159,g21179,g21244,g21253,g21261,g21269,g21501,g20522,g21536,
    g21540,g20542,g21572,g21576,g19067,g21605,g21609,g19084,g21634,g21774,
    g19121,g21787,II28305,g21788,g21789,g19128,II28318,g21799,g21800,g21801,
    II28323,g21802,g21803,g19135,g21806,II28330,g21807,g21808,g21809,II28335,
    g21810,g21811,g19138,g21813,II28341,g21814,g21815,g21816,II28346,g21817,
    g21819,II28351,g21820,g21821,g21823,II28365,g21844,II28369,g21846,II28374,
    g21849,II28380,g21856,g22175,g22190,g22199,g22205,g12451,g23319,g22385,
    g23688,g23742,g23797,g23850,g24239,g24244,g22317,g24245,g24252,g22342,
    g24254,g24257,g22365,g24258,g24965,g23922,g24978,g23954,g24989,g23983,
    g25000,g24013,g25183,g25186,g25190,g25195,g26320,g25852,g26367,g25873,
    g26410,g25885,g26451,g25890,g27738,g27743,g27751,g27756,II15167,II15168,
    II15169,g7855,II15183,II15184,II15185,g7875,II15190,II15191,II15192,g7876,
    II15204,II15205,II15206,g7895,II15211,II15212,II15213,g7896,II15237,
    II15238,II15239,g7922,II15244,II15245,II15246,g7923,II15276,II15277,
    II15278,g7970,II16879,II16880,II16881,g9883,II16965,II16966,II16967,g10003,
    II17059,II17060,II17061,g10095,II17149,II17150,II17151,g10185,II18106,
    II18107,II18108,g11188,II18113,II18114,II18115,g11189,II18190,II18191,
    II18192,g11262,II18197,II18198,II18199,g11263,II18204,II18205,II18206,
    g11264,II18280,II18281,II18282,g11330,II18287,II18288,II18289,g11331,
    II18368,II18369,II18370,g11410,II18799,II18800,II18801,g11621,II20031,
    II20032,II20033,g12988,II20048,II20049,II20050,g12999,II20429,II20430,
    II20431,g13348,II20465,II20466,II20467,g13370,II20504,II20505,II20506,
    g13399,II20743,II20744,II20745,g13507,g13893,g13915,g13934,g13957,g13971,
    g13990,g14027,g14041,g14060,g14118,g14132,g14233,g12780,g12819,g12857,
    g13401,g12898,g13286,g13313,g11622,g13332,g11643,g13375,g11660,II22062,
    II22063,II22064,g15814,g13024,g13310,g13331,g13353,g13354,g13374,g13404,
    II22282,II22283,II22284,II22316,II22317,II22318,II22630,g15978,II22631,
    II22632,II22705,g15661,II22706,II22707,II22884,II22885,II22886,II22900,
    II22901,II22902,II22917,II22918,II22919,II22924,II22925,II22926,II22936,
    II22937,II22938,II22945,II22946,II22947,II22952,II22953,II22954,II22962,
    II22963,II22964,II22972,II22973,II22974,II22981,II22982,II22983,II22988,
    II22989,II22990,II22998,II22999,II23000,II23008,II23009,II23010,II23018,
    II23019,II23020,II23027,II23028,II23029,II23034,II23035,II23036,II23045,
    II23046,II23047,II23055,II23056,II23057,II23065,II23066,II23067,II23074,
    II23075,II23076,II23082,II23083,II23084,II23093,II23094,II23095,II23103,
    II23104,II23105,II23113,II23114,II23115,II23123,II23124,II23125,II23131,
    II23132,II23133,II23142,II23143,II23144,II23152,II23153,II23154,II23161,
    II23162,II23163,II23171,II23172,II23173,II23179,II23180,II23181,II23190,
    II23191,II23192,II23198,II23199,II23200,II23207,II23208,II23209,II23217,
    II23218,II23219,II23225,II23226,II23227,II23233,II23234,II23235,II23242,
    II23243,II23244,II23256,II23257,II23258,II23264,II23265,II23266,II23277,
    II23278,II23279,II23806,II23807,II23808,II23878,II23879,II23880,II23893,
    II23894,II23895,II23941,II23942,II23943,II23958,II23959,II23960,II23966,
    II23967,II23968,II23981,II23982,II23983,II24005,II24006,II24007,II24015,
    II24016,II24017,II24028,II24029,II24030,II24036,II24037,II24038,II24053,
    II24054,II24055,II24061,II24062,II24063,II24076,II24077,II24078,II24091,
    II24092,II24093,II24102,II24103,II24104,II24110,II24111,II24112,II24123,
    II24124,II24125,II24131,II24132,II24133,II24148,II24149,II24150,II24156,
    II24157,II24158,II24178,II24179,II24180,II24186,II24187,II24188,II24194,
    II24195,II24196,II24205,II24206,II24207,II24213,II24214,II24215,II24226,
    II24227,II24228,II24234,II24235,II24236,II24251,II24252,II24253,II24263,
    II24264,II24265,II24271,II24272,II24273,II24278,II24279,II24280,II24290,
    II24291,II24292,II24298,II24299,II24300,II24306,II24307,II24308,II24317,
    II24318,II24319,II24325,II24326,II24327,II24338,II24339,II24340,II24351,
    II24352,II24353,II24361,II24362,II24363,II24372,II24373,II24374,II24380,
    II24381,II24382,II24387,II24388,II24389,II24399,II24400,II24401,II24407,
    II24408,II24409,II24415,II24416,II24417,II24426,II24427,II24428,II24436,
    II24437,II24438,II24443,II24444,II24445,II24452,II24453,II24454,II24464,
    II24465,II24466,II24474,II24475,II24476,II24485,II24486,II24487,II24493,
    II24494,II24495,II24500,II24501,II24502,II24512,II24513,II24514,II24520,
    II24521,II24522,II24530,II24531,II24532,II24537,II24538,II24539,II24544,
    II24545,II24546,II24553,II24554,II24555,II24565,II24566,II24567,II24575,
    II24576,II24577,II24586,II24587,II24588,II24594,II24595,II24596,II24601,
    II24602,II24603,II24611,II24612,II24613,II24624,II24625,II24626,II24632,
    II24633,II24634,II24639,II24640,II24641,II24646,II24647,II24648,II24655,
    II24656,II24657,II24667,II24668,II24669,II24677,II24678,II24679,II24694,
    II24695,II24696,II24702,II24703,II24704,II24709,II24710,II24711,II24716,
    II24717,II24718,II24725,II24726,II24727,II24743,II24744,II24745,II24751,
    II24752,II24753,II24763,II24764,II24765,II25030,II25031,II25032,II25532,
    II25533,II25534,II25539,II25540,II25541,II25560,II25561,II25562,II25571,
    II25572,II25573,II25578,II25579,II25580,II25595,II25596,II25597,II25605,
    II25606,II25607,II25616,II25617,II25618,II25623,II25624,II25625,II25633,
    II25634,II25635,II25643,II25644,II25645,II25653,II25654,II25655,II25664,
    II25665,II25666,II25671,II25672,II25673,II25681,II25682,II25683,II25690,
    II25691,II25692,II25700,II25701,II25702,II25710,II25711,II25712,II25721,
    II25722,II25723,II25731,II25732,II25733,II25740,II25741,II25742,II25750,
    II25751,II25752,II25761,II25762,II25763,II25771,II25772,II25773,II25781,
    II25782,II25783,II25790,II25791,II25792,II25800,II25801,II25802,II25809,
    II25810,II25811,II25819,II25820,II25821,II25829,II25830,II25831,II25838,
    II25839,II25840,II25846,II25847,II25848,II25855,II25856,II25857,II25865,
    II25866,II25867,II25880,II25881,II25882,II25888,II25889,II25890,II25897,
    II25898,II25899,II25913,II25914,II25915,II25921,II25922,II25923,II25938,
    II25939,II25940,g19219,II28189,II28190,II28191,g21660,II28217,II28218,
    II28219,g21689,II28247,II28248,II28249,g21725,II28271,II28272,II28273,
    g21751,g21848,g21850,g21855,g21857,g21858,g21859,g21860,g21862,g21863,
    g21864,g21865,g21866,g21868,g21869,g21870,g21871,g21873,g21874,g21875,
    g21877,g21879,g21881,g21885,g21888,g21048,g21065,II28726,g21887,II28727,
    II28728,II28741,g21890,II28742,II28743,II28753,g21893,II28754,II28755,
    II28765,g21901,II28766,II28767,g21211,g21219,g21230,g21235,g22809,g22844,
    g22846,g22850,g22879,g22881,g22885,g22914,g22916,g22920,g22939,g22941,
    g23066,g23051,g23080,g23070,g22999,g22174,g23096,g23083,g23013,g22189,
    g23113,g23099,g23029,g22198,g23046,g22204,g21980,g21975,g21987,g21981,
    g23135,g22288,g22000,g21988,g23376,g21968,g22308,g22013,g22001,g23387,
    g21971,g22336,g23394,g21973,g22361,g23402,II30790,II30791,II30792,II30868,
    II30869,II30870,II30952,II30953,II30954,II31035,II31036,II31037,g23906,
    g23936,g23937,g23938,g23953,g23968,g23969,g23970,g23973,g23982,g23997,
    g23998,g23999,g24002,g24003,g24012,g24027,g24028,g24034,g24036,g24037,
    g24046,g24052,g24054,g24056,g24057,g24058,g24065,g24067,g24069,g24070,
    g24071,g24078,g24080,g24081,g24082,g24089,g24090,g24091,g24093,II32265,
    II32266,II32267,II32284,II32285,II32286,II32295,II32296,II32297,II32308,
    II32309,II32310,II32323,II32324,II32325,II32333,II32334,II32335,II32345,
    II32346,II32347,II32355,II32356,II32357,II32368,II32369,II32370,II32378,
    II32379,II32380,II32391,II32392,II32393,II32400,II32401,II32402,II32409,
    II32410,II32411,II32422,II32423,II32424,II32430,II32431,II32432,II32443,
    II32444,II32445,II32451,II32452,II32453,II32460,II32461,II32462,II32468,
    II32469,II32470,II32478,II32479,II32480,II32490,II32491,II32492,II32498,
    II32499,II32500,II32509,II32510,II32511,II32518,II32519,II32520,II32526,
    II32527,II32528,II32538,II32539,II32540,II32546,II32547,II32548,II32559,
    II32560,II32561,II32567,II32568,II32569,II32575,II32576,II32577,II32586,
    II32587,II32588,II32595,II32596,II32597,II32607,II32608,II32609,II32615,
    II32616,II32617,II32624,II32625,II32626,II32633,II32634,II32635,II32645,
    II32646,II32647,II32659,II32660,II32661,II32668,II32669,II32670,II32677,
    g23823,II32678,II32679,II32686,II32687,II32688,II32695,g23858,II32696,
    II32697,II32708,g23892,II32709,II32710,II32724,g23913,II32725,II32726,
    g24517,g24530,g24543,g24555,II35020,II35021,II35022,g26859,II35034,II35035,
    II35036,g26865,II35042,II35043,II35044,g26867,II35057,II35058,II35059,
    g26874,g25699,g25569,g25631,g25772,g25648,g25708,g25826,g25725,g25781,
    g25861,g25798,g25835,II35123,g26107,g26096,II35124,II35125,II35701,II35702,
    II35703,g27379,II35714,II35715,II35716,g27382,g26989,g27012,g27038,g27066,
    II35904,g27051,II35905,II35906,II35944,g27078,II35945,II35946,II35974,
    g27094,II35975,II35976,II35992,g27106,II35993,II35994,g27415,g27436,g27455,
    g27471,II36256,g27527,II36257,II36258,g27801,II36270,g27549,II36271,
    II36272,g27809,II36289,g27565,II36290,II36291,g27830,II36300,II36301,
    II36302,II36314,g27575,II36315,II36316,g27846,II36591,g27529,II36592,
    II36593,II36666,g27551,II36667,II36668,II36731,g27567,II36732,II36733,
    II36779,g27577,II36780,II36781,II37295,II37296,II37297,g28384,II37303,
    II37304,II37305,g28386,II37311,II37312,II37313,g28388,II37322,II37323,
    II37324,g28391,II37356,g27824,g27811,II37357,II37358,II37813,II37814,
    II37815,g28842,II37822,II37823,II37824,g28845,II38378,II38379,II38380,
    II38810,g29303,II38811,II38812,II38820,g29313,II38821,II38822,II38831,
    g29324,II38832,II38833,II38841,g29333,II38842,II38843,II39323,II39324,
    II39325,g29911,II39331,II39332,II39333,g29913,II39339,II39340,II39341,
    g29915,II39347,II39348,II39349,g29917,II39359,g29766,II39360,II39361,
    g29923,II39367,g29767,II39368,II39369,g29925,II39375,g29768,II39376,
    II39377,g29927,II39384,g29718,g29710,II39385,II39386,II39391,g29769,
    II39392,II39393,g29931,II39532,II39533,II39534,g30034,II39539,II39540,
    II39541,g30035,II39689,II39690,II39691,II40558,II40559,II40560,g30768,
    II40571,II40572,II40573,g30771,II40587,II40588,II40589,g30775,II40603,
    II40604,II40605,g30779,II40627,g30602,g30594,II40628,II40629,II41010,
    II41011,II41012,g30926,II41017,II41018,II41019,g30927,II41064,II41065,
    II41066,g16020,g16036,g16058,g16082,g16094,g16120,g16171,g16230,g18352,
    g18430,g18447,g18503,g18520,g18567,g18584,g18617,g19160,g19165,g19171,
    g19177,g20878,g20895,g20914,g20938,g21083,g21618,g21646,g21677,g21706,
    g21738,g21762,g21778,g21793,g22144,g22165,g22181,g22186,g22195,g22210,
    g22216,g22227,g22985,g22987,g22990,g22997,g23009,g23025,g23042,g23061,
    g23386,g23393,g23401,g23408,g23427,g23433,g23461,g23477,g24227,g24234,
    g24242,g24249,g24428,g24486,g24490,g24492,g24493,g24497,g24500,g24502,
    g24503,g24506,g24509,g24512,g24514,g24515,g24516,g24520,g24523,g24526,
    g24528,g24533,g24536,g24546,g24558,g24566,g24575,g24613,g24622,g24624,
    g24637,g24638,g24656,g24657,g24675,g24708,g24717,g24720,g24728,g24731,
    g24736,g24739,g24742,g25076,g25077,g25078,g25081,g25082,g25085,g25091,
    g25099,g25125,g25127,g25129,g25208,g25216,g25226,g25238,g25273,g25311,
    g25426,g25962,g25967,g25974,g25979,g26042,g26044,g26046,g26049,g26050,
    g26055,g26081,g26084,g26090,g26103,g26140,g26560,g26583,g26607,g26630,
    g26799,g26800,g26801,g26802,g26873,g26882,g26891,g26901,g27175,g27179,
    g27184,g27188,g27250,g27251,g27252,g27254,g27478,g27501,g27521,g27546,
    g27629,g27631,g27655,g27658,g27736,g27742,g27747,g27755,g27869,g27886,
    g28185,g28189,g28191,g28192,g28654,g28656,g28658,g28661,g29126,g29127,
    g29128,g29129,g29399,g29403,g29406,g29409,g29736,g29744,g30618,g30625;

  dff DFF_0(CK,g2814,g16475);
  dff DFF_1(CK,g2817,g20571);
  dff DFF_2(CK,g2933,g20588);
  dff DFF_3(CK,g2950,g21951);
  dff DFF_4(CK,g2883,g23315);
  dff DFF_5(CK,g2888,g24423);
  dff DFF_6(CK,g2896,g25175);
  dff DFF_7(CK,g2892,g26019);
  dff DFF_8(CK,g2903,g26747);
  dff DFF_9(CK,g2900,g27237);
  dff DFF_10(CK,g2908,g27715);
  dff DFF_11(CK,g2912,g24424);
  dff DFF_12(CK,g2917,g25174);
  dff DFF_13(CK,g2924,g26020);
  dff DFF_14(CK,g2920,g26746);
  dff DFF_15(CK,g2984,g19061);
  dff DFF_16(CK,g2985,g19060);
  dff DFF_17(CK,g2930,g19062);
  dff DFF_18(CK,g2929,g2930);
  dff DFF_19(CK,g2879,g16494);
  dff DFF_20(CK,g2934,g16476);
  dff DFF_21(CK,g2935,g16477);
  dff DFF_22(CK,g2938,g16478);
  dff DFF_23(CK,g2941,g16479);
  dff DFF_24(CK,g2944,g16480);
  dff DFF_25(CK,g2947,g16481);
  dff DFF_26(CK,g2953,g16482);
  dff DFF_27(CK,g2956,g16483);
  dff DFF_28(CK,g2959,g16484);
  dff DFF_29(CK,g2962,g16485);
  dff DFF_30(CK,g2963,g16486);
  dff DFF_31(CK,g2966,g16487);
  dff DFF_32(CK,g2969,g16488);
  dff DFF_33(CK,g2972,g16489);
  dff DFF_34(CK,g2975,g16490);
  dff DFF_35(CK,g2978,g16491);
  dff DFF_36(CK,g2981,g16492);
  dff DFF_37(CK,g2874,g16493);
  dff DFF_38(CK,g1506,g20572);
  dff DFF_39(CK,g1501,g20573);
  dff DFF_40(CK,g1496,g20574);
  dff DFF_41(CK,g1491,g20575);
  dff DFF_42(CK,g1486,g20576);
  dff DFF_43(CK,g1481,g20577);
  dff DFF_44(CK,g1476,g20578);
  dff DFF_45(CK,g1471,g20579);
  dff DFF_46(CK,g2877,g23313);
  dff DFF_47(CK,g2861,g21960);
  dff DFF_48(CK,g813,g2861);
  dff DFF_49(CK,g2864,g21961);
  dff DFF_50(CK,g809,g2864);
  dff DFF_51(CK,g2867,g21962);
  dff DFF_52(CK,g805,g2867);
  dff DFF_53(CK,g2870,g21963);
  dff DFF_54(CK,g801,g2870);
  dff DFF_55(CK,g2818,g21947);
  dff DFF_56(CK,g797,g2818);
  dff DFF_57(CK,g2821,g21948);
  dff DFF_58(CK,g793,g2821);
  dff DFF_59(CK,g2824,g21949);
  dff DFF_60(CK,g789,g2824);
  dff DFF_61(CK,g2827,g21950);
  dff DFF_62(CK,g785,g2827);
  dff DFF_63(CK,g2830,g23312);
  dff DFF_64(CK,g2873,g2830);
  dff DFF_65(CK,g2833,g21952);
  dff DFF_66(CK,g125,g2833);
  dff DFF_67(CK,g2836,g21953);
  dff DFF_68(CK,g121,g2836);
  dff DFF_69(CK,g2839,g21954);
  dff DFF_70(CK,g117,g2839);
  dff DFF_71(CK,g2842,g21955);
  dff DFF_72(CK,g113,g2842);
  dff DFF_73(CK,g2845,g21956);
  dff DFF_74(CK,g109,g2845);
  dff DFF_75(CK,g2848,g21957);
  dff DFF_76(CK,g105,g2848);
  dff DFF_77(CK,g2851,g21958);
  dff DFF_78(CK,g101,g2851);
  dff DFF_79(CK,g2854,g21959);
  dff DFF_80(CK,g97,g2854);
  dff DFF_81(CK,g2858,g23316);
  dff DFF_82(CK,g2857,g2858);
  dff DFF_83(CK,g2200,g20587);
  dff DFF_84(CK,g2195,g20585);
  dff DFF_85(CK,g2190,g20586);
  dff DFF_86(CK,g2185,g20584);
  dff DFF_87(CK,g2180,g20583);
  dff DFF_88(CK,g2175,g20582);
  dff DFF_89(CK,g2170,g20581);
  dff DFF_90(CK,g2165,g20580);
  dff DFF_91(CK,g2878,g23314);
  dff DFF_92(CK,g3129,g13475);
  dff DFF_93(CK,g3117,g3129);
  dff DFF_94(CK,g3109,g3117);
  dff DFF_95(CK,g3210,g20630);
  dff DFF_96(CK,g3211,g20631);
  dff DFF_97(CK,g3084,g20632);
  dff DFF_98(CK,g3085,g20609);
  dff DFF_99(CK,g3086,g20610);
  dff DFF_100(CK,g3087,g20611);
  dff DFF_101(CK,g3091,g20612);
  dff DFF_102(CK,g3092,g20613);
  dff DFF_103(CK,g3093,g20614);
  dff DFF_104(CK,g3094,g20615);
  dff DFF_105(CK,g3095,g20616);
  dff DFF_106(CK,g3096,g20617);
  dff DFF_107(CK,g3097,g26751);
  dff DFF_108(CK,g3098,g26752);
  dff DFF_109(CK,g3099,g26753);
  dff DFF_110(CK,g3100,g29163);
  dff DFF_111(CK,g3101,g29164);
  dff DFF_112(CK,g3102,g29165);
  dff DFF_113(CK,g3103,g30120);
  dff DFF_114(CK,g3104,g30121);
  dff DFF_115(CK,g3105,g30122);
  dff DFF_116(CK,g3106,g30941);
  dff DFF_117(CK,g3107,g30942);
  dff DFF_118(CK,g3108,g30943);
  dff DFF_119(CK,g3155,g20618);
  dff DFF_120(CK,g3158,g20619);
  dff DFF_121(CK,g3161,g20620);
  dff DFF_122(CK,g3164,g20621);
  dff DFF_123(CK,g3167,g20622);
  dff DFF_124(CK,g3170,g20623);
  dff DFF_125(CK,g3173,g20624);
  dff DFF_126(CK,g3176,g20625);
  dff DFF_127(CK,g3179,g20626);
  dff DFF_128(CK,g3182,g20627);
  dff DFF_129(CK,g3185,g20628);
  dff DFF_130(CK,g3088,g20629);
  dff DFF_131(CK,g3191,g27717);
  dff DFF_132(CK,g3194,g28316);
  dff DFF_133(CK,g3197,g28317);
  dff DFF_134(CK,g3198,g28318);
  dff DFF_135(CK,g3201,g28704);
  dff DFF_136(CK,g3204,g28705);
  dff DFF_137(CK,g3207,g28706);
  dff DFF_138(CK,g3188,g29463);
  dff DFF_139(CK,g3133,g29656);
  dff DFF_140(CK,g3132,g28698);
  dff DFF_141(CK,g3128,g29166);
  dff DFF_142(CK,g3127,g28697);
  dff DFF_143(CK,g3126,g28315);
  dff DFF_144(CK,g3125,g28696);
  dff DFF_145(CK,g3124,g28314);
  dff DFF_146(CK,g3123,g28313);
  dff DFF_147(CK,g3120,g28695);
  dff DFF_148(CK,g3114,g28694);
  dff DFF_149(CK,g3113,g28693);
  dff DFF_150(CK,g3112,g28312);
  dff DFF_151(CK,g3110,g28311);
  dff DFF_152(CK,g3111,g28310);
  dff DFF_153(CK,g3139,g29461);
  dff DFF_154(CK,g3136,g28701);
  dff DFF_155(CK,g3134,g28700);
  dff DFF_156(CK,g3135,g28699);
  dff DFF_157(CK,g3151,g29462);
  dff DFF_158(CK,g3142,g28703);
  dff DFF_159(CK,g3147,g28702);
  dff DFF_160(CK,g185,g29657);
  dff DFF_161(CK,g138,g13405);
  dff DFF_162(CK,g135,g138);
  dff DFF_163(CK,g165,g135);
  dff DFF_164(CK,g130,g24259);
  dff DFF_165(CK,g131,g24260);
  dff DFF_166(CK,g129,g24261);
  dff DFF_167(CK,g133,g24262);
  dff DFF_168(CK,g134,g24263);
  dff DFF_169(CK,g132,g24264);
  dff DFF_170(CK,g142,g24265);
  dff DFF_171(CK,g143,g24266);
  dff DFF_172(CK,g141,g24267);
  dff DFF_173(CK,g145,g24268);
  dff DFF_174(CK,g146,g24269);
  dff DFF_175(CK,g144,g24270);
  dff DFF_176(CK,g148,g24271);
  dff DFF_177(CK,g149,g24272);
  dff DFF_178(CK,g147,g24273);
  dff DFF_179(CK,g151,g24274);
  dff DFF_180(CK,g152,g24275);
  dff DFF_181(CK,g150,g24276);
  dff DFF_182(CK,g154,g24277);
  dff DFF_183(CK,g155,g24278);
  dff DFF_184(CK,g153,g24279);
  dff DFF_185(CK,g157,g24280);
  dff DFF_186(CK,g158,g24281);
  dff DFF_187(CK,g156,g24282);
  dff DFF_188(CK,g160,g24283);
  dff DFF_189(CK,g161,g24284);
  dff DFF_190(CK,g159,g24285);
  dff DFF_191(CK,g163,g24286);
  dff DFF_192(CK,g164,g24287);
  dff DFF_193(CK,g162,g24288);
  dff DFF_194(CK,g169,g26679);
  dff DFF_195(CK,g170,g26680);
  dff DFF_196(CK,g168,g26681);
  dff DFF_197(CK,g172,g26682);
  dff DFF_198(CK,g173,g26683);
  dff DFF_199(CK,g171,g26684);
  dff DFF_200(CK,g175,g26685);
  dff DFF_201(CK,g176,g26686);
  dff DFF_202(CK,g174,g26687);
  dff DFF_203(CK,g178,g26688);
  dff DFF_204(CK,g179,g26689);
  dff DFF_205(CK,g177,g26690);
  dff DFF_206(CK,g186,g30506);
  dff DFF_207(CK,g189,g30507);
  dff DFF_208(CK,g192,g30508);
  dff DFF_209(CK,g231,g30842);
  dff DFF_210(CK,g234,g30843);
  dff DFF_211(CK,g237,g30844);
  dff DFF_212(CK,g195,g30836);
  dff DFF_213(CK,g198,g30837);
  dff DFF_214(CK,g201,g30838);
  dff DFF_215(CK,g240,g30845);
  dff DFF_216(CK,g243,g30846);
  dff DFF_217(CK,g246,g30847);
  dff DFF_218(CK,g204,g30509);
  dff DFF_219(CK,g207,g30510);
  dff DFF_220(CK,g210,g30511);
  dff DFF_221(CK,g249,g30515);
  dff DFF_222(CK,g252,g30516);
  dff DFF_223(CK,g255,g30517);
  dff DFF_224(CK,g213,g30512);
  dff DFF_225(CK,g216,g30513);
  dff DFF_226(CK,g219,g30514);
  dff DFF_227(CK,g258,g30518);
  dff DFF_228(CK,g261,g30519);
  dff DFF_229(CK,g264,g30520);
  dff DFF_230(CK,g222,g30839);
  dff DFF_231(CK,g225,g30840);
  dff DFF_232(CK,g228,g30841);
  dff DFF_233(CK,g267,g30848);
  dff DFF_234(CK,g270,g30849);
  dff DFF_235(CK,g273,g30850);
  dff DFF_236(CK,g92,g25983);
  dff DFF_237(CK,g88,g26678);
  dff DFF_238(CK,g83,g27189);
  dff DFF_239(CK,g79,g27683);
  dff DFF_240(CK,g74,g28206);
  dff DFF_241(CK,g70,g28673);
  dff DFF_242(CK,g65,g29131);
  dff DFF_243(CK,g61,g29413);
  dff DFF_244(CK,g56,g29627);
  dff DFF_245(CK,g52,g29794);
  dff DFF_246(CK,g180,g20555);
  dff DFF_247(CK,g182,g180);
  dff DFF_248(CK,g181,g182);
  dff DFF_249(CK,g276,g13406);
  dff DFF_250(CK,g405,g276);
  dff DFF_251(CK,g401,g405);
  dff DFF_252(CK,g309,g11496);
  dff DFF_253(CK,g354,g28207);
  dff DFF_254(CK,g343,g28208);
  dff DFF_255(CK,g346,g28209);
  dff DFF_256(CK,g369,g28210);
  dff DFF_257(CK,g358,g28211);
  dff DFF_258(CK,g361,g28212);
  dff DFF_259(CK,g384,g28213);
  dff DFF_260(CK,g373,g28214);
  dff DFF_261(CK,g376,g28215);
  dff DFF_262(CK,g398,g28216);
  dff DFF_263(CK,g388,g28217);
  dff DFF_264(CK,g391,g28218);
  dff DFF_265(CK,g408,g29414);
  dff DFF_266(CK,g411,g29415);
  dff DFF_267(CK,g414,g29416);
  dff DFF_268(CK,g417,g29631);
  dff DFF_269(CK,g420,g29632);
  dff DFF_270(CK,g423,g29633);
  dff DFF_271(CK,g427,g29417);
  dff DFF_272(CK,g428,g29418);
  dff DFF_273(CK,g426,g29419);
  dff DFF_274(CK,g429,g27684);
  dff DFF_275(CK,g432,g27685);
  dff DFF_276(CK,g435,g27686);
  dff DFF_277(CK,g438,g27687);
  dff DFF_278(CK,g441,g27688);
  dff DFF_279(CK,g444,g27689);
  dff DFF_280(CK,g448,g28674);
  dff DFF_281(CK,g449,g28675);
  dff DFF_282(CK,g447,g28676);
  dff DFF_283(CK,g312,g29795);
  dff DFF_284(CK,g313,g29796);
  dff DFF_285(CK,g314,g29797);
  dff DFF_286(CK,g315,g30851);
  dff DFF_287(CK,g316,g30852);
  dff DFF_288(CK,g317,g30853);
  dff DFF_289(CK,g318,g30710);
  dff DFF_290(CK,g319,g30711);
  dff DFF_291(CK,g320,g30712);
  dff DFF_292(CK,g322,g29628);
  dff DFF_293(CK,g323,g29629);
  dff DFF_294(CK,g321,g29630);
  dff DFF_295(CK,g403,g27191);
  dff DFF_296(CK,g404,g27192);
  dff DFF_297(CK,g402,g27193);
  dff DFF_298(CK,g450,g11509);
  dff DFF_299(CK,g451,g450);
  dff DFF_300(CK,g452,g11510);
  dff DFF_301(CK,g453,g452);
  dff DFF_302(CK,g454,g11511);
  dff DFF_303(CK,g279,g454);
  dff DFF_304(CK,g280,g11491);
  dff DFF_305(CK,g281,g280);
  dff DFF_306(CK,g282,g11492);
  dff DFF_307(CK,g283,g282);
  dff DFF_308(CK,g284,g11493);
  dff DFF_309(CK,g285,g284);
  dff DFF_310(CK,g286,g11494);
  dff DFF_311(CK,g287,g286);
  dff DFF_312(CK,g288,g11495);
  dff DFF_313(CK,g289,g288);
  dff DFF_314(CK,g290,g13407);
  dff DFF_315(CK,g291,g290);
  dff DFF_316(CK,g299,g19012);
  dff DFF_317(CK,g305,g23148);
  dff DFF_318(CK,g308,g23149);
  dff DFF_319(CK,g297,g23150);
  dff DFF_320(CK,g296,g23151);
  dff DFF_321(CK,g295,g23152);
  dff DFF_322(CK,g294,g23153);
  dff DFF_323(CK,g304,g19016);
  dff DFF_324(CK,g303,g19015);
  dff DFF_325(CK,g302,g19014);
  dff DFF_326(CK,g301,g19013);
  dff DFF_327(CK,g300,g25130);
  dff DFF_328(CK,g298,g27190);
  dff DFF_329(CK,g342,g11497);
  dff DFF_330(CK,g349,g342);
  dff DFF_331(CK,g350,g11498);
  dff DFF_332(CK,g351,g350);
  dff DFF_333(CK,g352,g11499);
  dff DFF_334(CK,g353,g352);
  dff DFF_335(CK,g357,g11500);
  dff DFF_336(CK,g364,g357);
  dff DFF_337(CK,g365,g11501);
  dff DFF_338(CK,g366,g365);
  dff DFF_339(CK,g367,g11502);
  dff DFF_340(CK,g368,g367);
  dff DFF_341(CK,g372,g11503);
  dff DFF_342(CK,g379,g372);
  dff DFF_343(CK,g380,g11504);
  dff DFF_344(CK,g381,g380);
  dff DFF_345(CK,g382,g11505);
  dff DFF_346(CK,g383,g382);
  dff DFF_347(CK,g387,g11506);
  dff DFF_348(CK,g394,g387);
  dff DFF_349(CK,g395,g11507);
  dff DFF_350(CK,g396,g395);
  dff DFF_351(CK,g397,g11508);
  dff DFF_352(CK,g324,g397);
  dff DFF_353(CK,g325,g13408);
  dff DFF_354(CK,g331,g325);
  dff DFF_355(CK,g337,g331);
  dff DFF_356(CK,g545,g13419);
  dff DFF_357(CK,g551,g545);
  dff DFF_358(CK,g550,g551);
  dff DFF_359(CK,g554,g23160);
  dff DFF_360(CK,g557,g20556);
  dff DFF_361(CK,g510,g20557);
  dff DFF_362(CK,g513,g16467);
  dff DFF_363(CK,g523,g513);
  dff DFF_364(CK,g524,g523);
  dff DFF_365(CK,g564,g11512);
  dff DFF_366(CK,g569,g564);
  dff DFF_367(CK,g570,g11515);
  dff DFF_368(CK,g571,g570);
  dff DFF_369(CK,g572,g11516);
  dff DFF_370(CK,g573,g572);
  dff DFF_371(CK,g574,g11517);
  dff DFF_372(CK,g565,g574);
  dff DFF_373(CK,g566,g11513);
  dff DFF_374(CK,g567,g566);
  dff DFF_375(CK,g568,g11514);
  dff DFF_376(CK,g489,g568);
  dff DFF_377(CK,g474,g13409);
  dff DFF_378(CK,g481,g474);
  dff DFF_379(CK,g485,g481);
  dff DFF_380(CK,g486,g24292);
  dff DFF_381(CK,g487,g24293);
  dff DFF_382(CK,g488,g24294);
  dff DFF_383(CK,g455,g25139);
  dff DFF_384(CK,g458,g25131);
  dff DFF_385(CK,g461,g25132);
  dff DFF_386(CK,g477,g25136);
  dff DFF_387(CK,g478,g25137);
  dff DFF_388(CK,g479,g25138);
  dff DFF_389(CK,g480,g24289);
  dff DFF_390(CK,g484,g24290);
  dff DFF_391(CK,g464,g24291);
  dff DFF_392(CK,g465,g25133);
  dff DFF_393(CK,g468,g25134);
  dff DFF_394(CK,g471,g25135);
  dff DFF_395(CK,g528,g16468);
  dff DFF_396(CK,g535,g528);
  dff DFF_397(CK,g542,g535);
  dff DFF_398(CK,g543,g19021);
  dff DFF_399(CK,g544,g543);
  dff DFF_400(CK,g548,g23159);
  dff DFF_401(CK,g549,g19022);
  dff DFF_402(CK,g499,g549);
  dff DFF_403(CK,g558,g19023);
  dff DFF_404(CK,g559,g558);
  dff DFF_405(CK,g576,g28219);
  dff DFF_406(CK,g577,g28220);
  dff DFF_407(CK,g575,g28221);
  dff DFF_408(CK,g579,g28222);
  dff DFF_409(CK,g580,g28223);
  dff DFF_410(CK,g578,g28224);
  dff DFF_411(CK,g582,g28225);
  dff DFF_412(CK,g583,g28226);
  dff DFF_413(CK,g581,g28227);
  dff DFF_414(CK,g585,g28228);
  dff DFF_415(CK,g586,g28229);
  dff DFF_416(CK,g584,g28230);
  dff DFF_417(CK,g587,g25985);
  dff DFF_418(CK,g590,g25986);
  dff DFF_419(CK,g593,g25987);
  dff DFF_420(CK,g596,g25988);
  dff DFF_421(CK,g599,g25989);
  dff DFF_422(CK,g602,g25990);
  dff DFF_423(CK,g614,g29135);
  dff DFF_424(CK,g617,g29136);
  dff DFF_425(CK,g620,g29137);
  dff DFF_426(CK,g605,g29132);
  dff DFF_427(CK,g608,g29133);
  dff DFF_428(CK,g611,g29134);
  dff DFF_429(CK,g490,g27194);
  dff DFF_430(CK,g493,g27195);
  dff DFF_431(CK,g496,g27196);
  dff DFF_432(CK,g506,g8284);
  dff DFF_433(CK,g507,g24295);
  dff DFF_434(CK,g508,g19017);
  dff DFF_435(CK,g509,g19018);
  dff DFF_436(CK,g514,g19019);
  dff DFF_437(CK,g515,g19020);
  dff DFF_438(CK,g516,g23158);
  dff DFF_439(CK,g517,g23157);
  dff DFF_440(CK,g518,g23156);
  dff DFF_441(CK,g519,g23155);
  dff DFF_442(CK,g520,g23154);
  dff DFF_443(CK,g525,g520);
  dff DFF_444(CK,g529,g13410);
  dff DFF_445(CK,g530,g13411);
  dff DFF_446(CK,g531,g13412);
  dff DFF_447(CK,g532,g13413);
  dff DFF_448(CK,g533,g13414);
  dff DFF_449(CK,g534,g13415);
  dff DFF_450(CK,g536,g13416);
  dff DFF_451(CK,g537,g13417);
  dff DFF_452(CK,g538,g25984);
  dff DFF_453(CK,g541,g13418);
  dff DFF_454(CK,g623,g13420);
  dff DFF_455(CK,g626,g623);
  dff DFF_456(CK,g629,g626);
  dff DFF_457(CK,g630,g20558);
  dff DFF_458(CK,g659,g21943);
  dff DFF_459(CK,g640,g23161);
  dff DFF_460(CK,g633,g24296);
  dff DFF_461(CK,g653,g25140);
  dff DFF_462(CK,g646,g25991);
  dff DFF_463(CK,g660,g26691);
  dff DFF_464(CK,g672,g27197);
  dff DFF_465(CK,g666,g27690);
  dff DFF_466(CK,g679,g28231);
  dff DFF_467(CK,g686,g28677);
  dff DFF_468(CK,g692,g29138);
  dff DFF_469(CK,g699,g23162);
  dff DFF_470(CK,g700,g23163);
  dff DFF_471(CK,g698,g23164);
  dff DFF_472(CK,g702,g23165);
  dff DFF_473(CK,g703,g23166);
  dff DFF_474(CK,g701,g23167);
  dff DFF_475(CK,g705,g23168);
  dff DFF_476(CK,g706,g23169);
  dff DFF_477(CK,g704,g23170);
  dff DFF_478(CK,g708,g23171);
  dff DFF_479(CK,g709,g23172);
  dff DFF_480(CK,g707,g23173);
  dff DFF_481(CK,g711,g23174);
  dff DFF_482(CK,g712,g23175);
  dff DFF_483(CK,g710,g23176);
  dff DFF_484(CK,g714,g23177);
  dff DFF_485(CK,g715,g23178);
  dff DFF_486(CK,g713,g23179);
  dff DFF_487(CK,g717,g23180);
  dff DFF_488(CK,g718,g23181);
  dff DFF_489(CK,g716,g23182);
  dff DFF_490(CK,g720,g23183);
  dff DFF_491(CK,g721,g23184);
  dff DFF_492(CK,g719,g23185);
  dff DFF_493(CK,g723,g23186);
  dff DFF_494(CK,g724,g23187);
  dff DFF_495(CK,g722,g23188);
  dff DFF_496(CK,g726,g23189);
  dff DFF_497(CK,g727,g23190);
  dff DFF_498(CK,g725,g23191);
  dff DFF_499(CK,g729,g23192);
  dff DFF_500(CK,g730,g23193);
  dff DFF_501(CK,g728,g23194);
  dff DFF_502(CK,g732,g23195);
  dff DFF_503(CK,g733,g23196);
  dff DFF_504(CK,g731,g23197);
  dff DFF_505(CK,g735,g26692);
  dff DFF_506(CK,g736,g26693);
  dff DFF_507(CK,g734,g26694);
  dff DFF_508(CK,g738,g24297);
  dff DFF_509(CK,g739,g24298);
  dff DFF_510(CK,g737,g24299);
  dff DFF_511(CK,g826,g13421);
  dff DFF_512(CK,g823,g826);
  dff DFF_513(CK,g853,g823);
  dff DFF_514(CK,g818,g24300);
  dff DFF_515(CK,g819,g24301);
  dff DFF_516(CK,g817,g24302);
  dff DFF_517(CK,g821,g24303);
  dff DFF_518(CK,g822,g24304);
  dff DFF_519(CK,g820,g24305);
  dff DFF_520(CK,g830,g24306);
  dff DFF_521(CK,g831,g24307);
  dff DFF_522(CK,g829,g24308);
  dff DFF_523(CK,g833,g24309);
  dff DFF_524(CK,g834,g24310);
  dff DFF_525(CK,g832,g24311);
  dff DFF_526(CK,g836,g24312);
  dff DFF_527(CK,g837,g24313);
  dff DFF_528(CK,g835,g24314);
  dff DFF_529(CK,g839,g24315);
  dff DFF_530(CK,g840,g24316);
  dff DFF_531(CK,g838,g24317);
  dff DFF_532(CK,g842,g24318);
  dff DFF_533(CK,g843,g24319);
  dff DFF_534(CK,g841,g24320);
  dff DFF_535(CK,g845,g24321);
  dff DFF_536(CK,g846,g24322);
  dff DFF_537(CK,g844,g24323);
  dff DFF_538(CK,g848,g24324);
  dff DFF_539(CK,g849,g24325);
  dff DFF_540(CK,g847,g24326);
  dff DFF_541(CK,g851,g24327);
  dff DFF_542(CK,g852,g24328);
  dff DFF_543(CK,g850,g24329);
  dff DFF_544(CK,g857,g26696);
  dff DFF_545(CK,g858,g26697);
  dff DFF_546(CK,g856,g26698);
  dff DFF_547(CK,g860,g26699);
  dff DFF_548(CK,g861,g26700);
  dff DFF_549(CK,g859,g26701);
  dff DFF_550(CK,g863,g26702);
  dff DFF_551(CK,g864,g26703);
  dff DFF_552(CK,g862,g26704);
  dff DFF_553(CK,g866,g26705);
  dff DFF_554(CK,g867,g26706);
  dff DFF_555(CK,g865,g26707);
  dff DFF_556(CK,g873,g30521);
  dff DFF_557(CK,g876,g30522);
  dff DFF_558(CK,g879,g30523);
  dff DFF_559(CK,g918,g30860);
  dff DFF_560(CK,g921,g30861);
  dff DFF_561(CK,g924,g30862);
  dff DFF_562(CK,g882,g30854);
  dff DFF_563(CK,g885,g30855);
  dff DFF_564(CK,g888,g30856);
  dff DFF_565(CK,g927,g30863);
  dff DFF_566(CK,g930,g30864);
  dff DFF_567(CK,g933,g30865);
  dff DFF_568(CK,g891,g30524);
  dff DFF_569(CK,g894,g30525);
  dff DFF_570(CK,g897,g30526);
  dff DFF_571(CK,g936,g30530);
  dff DFF_572(CK,g939,g30531);
  dff DFF_573(CK,g942,g30532);
  dff DFF_574(CK,g900,g30527);
  dff DFF_575(CK,g903,g30528);
  dff DFF_576(CK,g906,g30529);
  dff DFF_577(CK,g945,g30533);
  dff DFF_578(CK,g948,g30534);
  dff DFF_579(CK,g951,g30535);
  dff DFF_580(CK,g909,g30857);
  dff DFF_581(CK,g912,g30858);
  dff DFF_582(CK,g915,g30859);
  dff DFF_583(CK,g954,g30866);
  dff DFF_584(CK,g957,g30867);
  dff DFF_585(CK,g960,g30868);
  dff DFF_586(CK,g780,g25992);
  dff DFF_587(CK,g776,g26695);
  dff DFF_588(CK,g771,g27198);
  dff DFF_589(CK,g767,g27691);
  dff DFF_590(CK,g762,g28232);
  dff DFF_591(CK,g758,g28678);
  dff DFF_592(CK,g753,g29139);
  dff DFF_593(CK,g749,g29420);
  dff DFF_594(CK,g744,g29634);
  dff DFF_595(CK,g740,g29798);
  dff DFF_596(CK,g868,g20559);
  dff DFF_597(CK,g870,g868);
  dff DFF_598(CK,g869,g870);
  dff DFF_599(CK,g963,g13422);
  dff DFF_600(CK,g1092,g963);
  dff DFF_601(CK,g1088,g1092);
  dff DFF_602(CK,g996,g11523);
  dff DFF_603(CK,g1041,g28233);
  dff DFF_604(CK,g1030,g28234);
  dff DFF_605(CK,g1033,g28235);
  dff DFF_606(CK,g1056,g28236);
  dff DFF_607(CK,g1045,g28237);
  dff DFF_608(CK,g1048,g28238);
  dff DFF_609(CK,g1071,g28239);
  dff DFF_610(CK,g1060,g28240);
  dff DFF_611(CK,g1063,g28241);
  dff DFF_612(CK,g1085,g28242);
  dff DFF_613(CK,g1075,g28243);
  dff DFF_614(CK,g1078,g28244);
  dff DFF_615(CK,g1095,g29421);
  dff DFF_616(CK,g1098,g29422);
  dff DFF_617(CK,g1101,g29423);
  dff DFF_618(CK,g1104,g29638);
  dff DFF_619(CK,g1107,g29639);
  dff DFF_620(CK,g1110,g29640);
  dff DFF_621(CK,g1114,g29424);
  dff DFF_622(CK,g1115,g29425);
  dff DFF_623(CK,g1113,g29426);
  dff DFF_624(CK,g1116,g27692);
  dff DFF_625(CK,g1119,g27693);
  dff DFF_626(CK,g1122,g27694);
  dff DFF_627(CK,g1125,g27695);
  dff DFF_628(CK,g1128,g27696);
  dff DFF_629(CK,g1131,g27697);
  dff DFF_630(CK,g1135,g28679);
  dff DFF_631(CK,g1136,g28680);
  dff DFF_632(CK,g1134,g28681);
  dff DFF_633(CK,g999,g29799);
  dff DFF_634(CK,g1000,g29800);
  dff DFF_635(CK,g1001,g29801);
  dff DFF_636(CK,g1002,g30869);
  dff DFF_637(CK,g1003,g30870);
  dff DFF_638(CK,g1004,g30871);
  dff DFF_639(CK,g1005,g30713);
  dff DFF_640(CK,g1006,g30714);
  dff DFF_641(CK,g1007,g30715);
  dff DFF_642(CK,g1009,g29635);
  dff DFF_643(CK,g1010,g29636);
  dff DFF_644(CK,g1008,g29637);
  dff DFF_645(CK,g1090,g27206);
  dff DFF_646(CK,g1091,g27207);
  dff DFF_647(CK,g1089,g27208);
  dff DFF_648(CK,g1137,g11536);
  dff DFF_649(CK,g1138,g1137);
  dff DFF_650(CK,g1139,g11537);
  dff DFF_651(CK,g1140,g1139);
  dff DFF_652(CK,g1141,g11538);
  dff DFF_653(CK,g966,g1141);
  dff DFF_654(CK,g967,g11518);
  dff DFF_655(CK,g968,g967);
  dff DFF_656(CK,g969,g11519);
  dff DFF_657(CK,g970,g969);
  dff DFF_658(CK,g971,g11520);
  dff DFF_659(CK,g972,g971);
  dff DFF_660(CK,g973,g11521);
  dff DFF_661(CK,g974,g973);
  dff DFF_662(CK,g975,g11522);
  dff DFF_663(CK,g976,g975);
  dff DFF_664(CK,g977,g13423);
  dff DFF_665(CK,g978,g977);
  dff DFF_666(CK,g986,g19024);
  dff DFF_667(CK,g992,g27200);
  dff DFF_668(CK,g995,g27201);
  dff DFF_669(CK,g984,g27202);
  dff DFF_670(CK,g983,g27203);
  dff DFF_671(CK,g982,g27204);
  dff DFF_672(CK,g981,g27205);
  dff DFF_673(CK,g991,g19028);
  dff DFF_674(CK,g990,g19027);
  dff DFF_675(CK,g989,g19026);
  dff DFF_676(CK,g988,g19025);
  dff DFF_677(CK,g987,g25141);
  dff DFF_678(CK,g985,g27199);
  dff DFF_679(CK,g1029,g11524);
  dff DFF_680(CK,g1036,g1029);
  dff DFF_681(CK,g1037,g11525);
  dff DFF_682(CK,g1038,g1037);
  dff DFF_683(CK,g1039,g11526);
  dff DFF_684(CK,g1040,g1039);
  dff DFF_685(CK,g1044,g11527);
  dff DFF_686(CK,g1051,g1044);
  dff DFF_687(CK,g1052,g11528);
  dff DFF_688(CK,g1053,g1052);
  dff DFF_689(CK,g1054,g11529);
  dff DFF_690(CK,g1055,g1054);
  dff DFF_691(CK,g1059,g11530);
  dff DFF_692(CK,g1066,g1059);
  dff DFF_693(CK,g1067,g11531);
  dff DFF_694(CK,g1068,g1067);
  dff DFF_695(CK,g1069,g11532);
  dff DFF_696(CK,g1070,g1069);
  dff DFF_697(CK,g1074,g11533);
  dff DFF_698(CK,g1081,g1074);
  dff DFF_699(CK,g1082,g11534);
  dff DFF_700(CK,g1083,g1082);
  dff DFF_701(CK,g1084,g11535);
  dff DFF_702(CK,g1011,g1084);
  dff DFF_703(CK,g1012,g13424);
  dff DFF_704(CK,g1018,g1012);
  dff DFF_705(CK,g1024,g1018);
  dff DFF_706(CK,g1231,g13435);
  dff DFF_707(CK,g1237,g1231);
  dff DFF_708(CK,g1236,g1237);
  dff DFF_709(CK,g1240,g23198);
  dff DFF_710(CK,g1243,g20560);
  dff DFF_711(CK,g1196,g20561);
  dff DFF_712(CK,g1199,g16469);
  dff DFF_713(CK,g1209,g1199);
  dff DFF_714(CK,g1210,g1209);
  dff DFF_715(CK,g1250,g11539);
  dff DFF_716(CK,g1255,g1250);
  dff DFF_717(CK,g1256,g11542);
  dff DFF_718(CK,g1257,g1256);
  dff DFF_719(CK,g1258,g11543);
  dff DFF_720(CK,g1259,g1258);
  dff DFF_721(CK,g1260,g11544);
  dff DFF_722(CK,g1251,g1260);
  dff DFF_723(CK,g1252,g11540);
  dff DFF_724(CK,g1253,g1252);
  dff DFF_725(CK,g1254,g11541);
  dff DFF_726(CK,g1176,g1254);
  dff DFF_727(CK,g1161,g13425);
  dff DFF_728(CK,g1168,g1161);
  dff DFF_729(CK,g1172,g1168);
  dff DFF_730(CK,g1173,g24333);
  dff DFF_731(CK,g1174,g24334);
  dff DFF_732(CK,g1175,g24335);
  dff DFF_733(CK,g1142,g25150);
  dff DFF_734(CK,g1145,g25142);
  dff DFF_735(CK,g1148,g25143);
  dff DFF_736(CK,g1164,g25147);
  dff DFF_737(CK,g1165,g25148);
  dff DFF_738(CK,g1166,g25149);
  dff DFF_739(CK,g1167,g24330);
  dff DFF_740(CK,g1171,g24331);
  dff DFF_741(CK,g1151,g24332);
  dff DFF_742(CK,g1152,g25144);
  dff DFF_743(CK,g1155,g25145);
  dff DFF_744(CK,g1158,g25146);
  dff DFF_745(CK,g1214,g16470);
  dff DFF_746(CK,g1221,g1214);
  dff DFF_747(CK,g1228,g1221);
  dff DFF_748(CK,g1229,g19033);
  dff DFF_749(CK,g1230,g1229);
  dff DFF_750(CK,g1234,g27217);
  dff DFF_751(CK,g1235,g19034);
  dff DFF_752(CK,g1186,g1235);
  dff DFF_753(CK,g1244,g19035);
  dff DFF_754(CK,g1245,g1244);
  dff DFF_755(CK,g1262,g28245);
  dff DFF_756(CK,g1263,g28246);
  dff DFF_757(CK,g1261,g28247);
  dff DFF_758(CK,g1265,g28248);
  dff DFF_759(CK,g1266,g28249);
  dff DFF_760(CK,g1264,g28250);
  dff DFF_761(CK,g1268,g28251);
  dff DFF_762(CK,g1269,g28252);
  dff DFF_763(CK,g1267,g28253);
  dff DFF_764(CK,g1271,g28254);
  dff DFF_765(CK,g1272,g28255);
  dff DFF_766(CK,g1270,g28256);
  dff DFF_767(CK,g1273,g25994);
  dff DFF_768(CK,g1276,g25995);
  dff DFF_769(CK,g1279,g25996);
  dff DFF_770(CK,g1282,g25997);
  dff DFF_771(CK,g1285,g25998);
  dff DFF_772(CK,g1288,g25999);
  dff DFF_773(CK,g1300,g29143);
  dff DFF_774(CK,g1303,g29144);
  dff DFF_775(CK,g1306,g29145);
  dff DFF_776(CK,g1291,g29140);
  dff DFF_777(CK,g1294,g29141);
  dff DFF_778(CK,g1297,g29142);
  dff DFF_779(CK,g1177,g27209);
  dff DFF_780(CK,g1180,g27210);
  dff DFF_781(CK,g1183,g27211);
  dff DFF_782(CK,g1192,g8293);
  dff DFF_783(CK,g1193,g24336);
  dff DFF_784(CK,g1194,g19029);
  dff DFF_785(CK,g1195,g19030);
  dff DFF_786(CK,g1200,g19031);
  dff DFF_787(CK,g1201,g19032);
  dff DFF_788(CK,g1202,g27216);
  dff DFF_789(CK,g1203,g27215);
  dff DFF_790(CK,g1204,g27214);
  dff DFF_791(CK,g1205,g27213);
  dff DFF_792(CK,g1206,g27212);
  dff DFF_793(CK,g1211,g1206);
  dff DFF_794(CK,g1215,g13426);
  dff DFF_795(CK,g1216,g13427);
  dff DFF_796(CK,g1217,g13428);
  dff DFF_797(CK,g1218,g13429);
  dff DFF_798(CK,g1219,g13430);
  dff DFF_799(CK,g1220,g13431);
  dff DFF_800(CK,g1222,g13432);
  dff DFF_801(CK,g1223,g13433);
  dff DFF_802(CK,g1224,g25993);
  dff DFF_803(CK,g1227,g13434);
  dff DFF_804(CK,g1309,g13436);
  dff DFF_805(CK,g1312,g1309);
  dff DFF_806(CK,g1315,g1312);
  dff DFF_807(CK,g1316,g20562);
  dff DFF_808(CK,g1345,g21944);
  dff DFF_809(CK,g1326,g23199);
  dff DFF_810(CK,g1319,g24337);
  dff DFF_811(CK,g1339,g25151);
  dff DFF_812(CK,g1332,g26000);
  dff DFF_813(CK,g1346,g26708);
  dff DFF_814(CK,g1358,g27218);
  dff DFF_815(CK,g1352,g27698);
  dff DFF_816(CK,g1365,g28257);
  dff DFF_817(CK,g1372,g28682);
  dff DFF_818(CK,g1378,g29146);
  dff DFF_819(CK,g1385,g23200);
  dff DFF_820(CK,g1386,g23201);
  dff DFF_821(CK,g1384,g23202);
  dff DFF_822(CK,g1388,g23203);
  dff DFF_823(CK,g1389,g23204);
  dff DFF_824(CK,g1387,g23205);
  dff DFF_825(CK,g1391,g23206);
  dff DFF_826(CK,g1392,g23207);
  dff DFF_827(CK,g1390,g23208);
  dff DFF_828(CK,g1394,g23209);
  dff DFF_829(CK,g1395,g23210);
  dff DFF_830(CK,g1393,g23211);
  dff DFF_831(CK,g1397,g23212);
  dff DFF_832(CK,g1398,g23213);
  dff DFF_833(CK,g1396,g23214);
  dff DFF_834(CK,g1400,g23215);
  dff DFF_835(CK,g1401,g23216);
  dff DFF_836(CK,g1399,g23217);
  dff DFF_837(CK,g1403,g23218);
  dff DFF_838(CK,g1404,g23219);
  dff DFF_839(CK,g1402,g23220);
  dff DFF_840(CK,g1406,g23221);
  dff DFF_841(CK,g1407,g23222);
  dff DFF_842(CK,g1405,g23223);
  dff DFF_843(CK,g1409,g23224);
  dff DFF_844(CK,g1410,g23225);
  dff DFF_845(CK,g1408,g23226);
  dff DFF_846(CK,g1412,g23227);
  dff DFF_847(CK,g1413,g23228);
  dff DFF_848(CK,g1411,g23229);
  dff DFF_849(CK,g1415,g23230);
  dff DFF_850(CK,g1416,g23231);
  dff DFF_851(CK,g1414,g23232);
  dff DFF_852(CK,g1418,g23233);
  dff DFF_853(CK,g1419,g23234);
  dff DFF_854(CK,g1417,g23235);
  dff DFF_855(CK,g1421,g26709);
  dff DFF_856(CK,g1422,g26710);
  dff DFF_857(CK,g1420,g26711);
  dff DFF_858(CK,g1424,g24338);
  dff DFF_859(CK,g1425,g24339);
  dff DFF_860(CK,g1423,g24340);
  dff DFF_861(CK,g1520,g13437);
  dff DFF_862(CK,g1517,g1520);
  dff DFF_863(CK,g1547,g1517);
  dff DFF_864(CK,g1512,g24341);
  dff DFF_865(CK,g1513,g24342);
  dff DFF_866(CK,g1511,g24343);
  dff DFF_867(CK,g1515,g24344);
  dff DFF_868(CK,g1516,g24345);
  dff DFF_869(CK,g1514,g24346);
  dff DFF_870(CK,g1524,g24347);
  dff DFF_871(CK,g1525,g24348);
  dff DFF_872(CK,g1523,g24349);
  dff DFF_873(CK,g1527,g24350);
  dff DFF_874(CK,g1528,g24351);
  dff DFF_875(CK,g1526,g24352);
  dff DFF_876(CK,g1530,g24353);
  dff DFF_877(CK,g1531,g24354);
  dff DFF_878(CK,g1529,g24355);
  dff DFF_879(CK,g1533,g24356);
  dff DFF_880(CK,g1534,g24357);
  dff DFF_881(CK,g1532,g24358);
  dff DFF_882(CK,g1536,g24359);
  dff DFF_883(CK,g1537,g24360);
  dff DFF_884(CK,g1535,g24361);
  dff DFF_885(CK,g1539,g24362);
  dff DFF_886(CK,g1540,g24363);
  dff DFF_887(CK,g1538,g24364);
  dff DFF_888(CK,g1542,g24365);
  dff DFF_889(CK,g1543,g24366);
  dff DFF_890(CK,g1541,g24367);
  dff DFF_891(CK,g1545,g24368);
  dff DFF_892(CK,g1546,g24369);
  dff DFF_893(CK,g1544,g24370);
  dff DFF_894(CK,g1551,g26713);
  dff DFF_895(CK,g1552,g26714);
  dff DFF_896(CK,g1550,g26715);
  dff DFF_897(CK,g1554,g26716);
  dff DFF_898(CK,g1555,g26717);
  dff DFF_899(CK,g1553,g26718);
  dff DFF_900(CK,g1557,g26719);
  dff DFF_901(CK,g1558,g26720);
  dff DFF_902(CK,g1556,g26721);
  dff DFF_903(CK,g1560,g26722);
  dff DFF_904(CK,g1561,g26723);
  dff DFF_905(CK,g1559,g26724);
  dff DFF_906(CK,g1567,g30536);
  dff DFF_907(CK,g1570,g30537);
  dff DFF_908(CK,g1573,g30538);
  dff DFF_909(CK,g1612,g30878);
  dff DFF_910(CK,g1615,g30879);
  dff DFF_911(CK,g1618,g30880);
  dff DFF_912(CK,g1576,g30872);
  dff DFF_913(CK,g1579,g30873);
  dff DFF_914(CK,g1582,g30874);
  dff DFF_915(CK,g1621,g30881);
  dff DFF_916(CK,g1624,g30882);
  dff DFF_917(CK,g1627,g30883);
  dff DFF_918(CK,g1585,g30539);
  dff DFF_919(CK,g1588,g30540);
  dff DFF_920(CK,g1591,g30541);
  dff DFF_921(CK,g1630,g30545);
  dff DFF_922(CK,g1633,g30546);
  dff DFF_923(CK,g1636,g30547);
  dff DFF_924(CK,g1594,g30542);
  dff DFF_925(CK,g1597,g30543);
  dff DFF_926(CK,g1600,g30544);
  dff DFF_927(CK,g1639,g30548);
  dff DFF_928(CK,g1642,g30549);
  dff DFF_929(CK,g1645,g30550);
  dff DFF_930(CK,g1603,g30875);
  dff DFF_931(CK,g1606,g30876);
  dff DFF_932(CK,g1609,g30877);
  dff DFF_933(CK,g1648,g30884);
  dff DFF_934(CK,g1651,g30885);
  dff DFF_935(CK,g1654,g30886);
  dff DFF_936(CK,g1466,g26001);
  dff DFF_937(CK,g1462,g26712);
  dff DFF_938(CK,g1457,g27219);
  dff DFF_939(CK,g1453,g27699);
  dff DFF_940(CK,g1448,g28258);
  dff DFF_941(CK,g1444,g28683);
  dff DFF_942(CK,g1439,g29147);
  dff DFF_943(CK,g1435,g29427);
  dff DFF_944(CK,g1430,g29641);
  dff DFF_945(CK,g1426,g29802);
  dff DFF_946(CK,g1562,g20563);
  dff DFF_947(CK,g1564,g1562);
  dff DFF_948(CK,g1563,g1564);
  dff DFF_949(CK,g1657,g13438);
  dff DFF_950(CK,g1786,g1657);
  dff DFF_951(CK,g1782,g1786);
  dff DFF_952(CK,g1690,g11550);
  dff DFF_953(CK,g1735,g28259);
  dff DFF_954(CK,g1724,g28260);
  dff DFF_955(CK,g1727,g28261);
  dff DFF_956(CK,g1750,g28262);
  dff DFF_957(CK,g1739,g28263);
  dff DFF_958(CK,g1742,g28264);
  dff DFF_959(CK,g1765,g28265);
  dff DFF_960(CK,g1754,g28266);
  dff DFF_961(CK,g1757,g28267);
  dff DFF_962(CK,g1779,g28268);
  dff DFF_963(CK,g1769,g28269);
  dff DFF_964(CK,g1772,g28270);
  dff DFF_965(CK,g1789,g29434);
  dff DFF_966(CK,g1792,g29435);
  dff DFF_967(CK,g1795,g29436);
  dff DFF_968(CK,g1798,g29645);
  dff DFF_969(CK,g1801,g29646);
  dff DFF_970(CK,g1804,g29647);
  dff DFF_971(CK,g1808,g29437);
  dff DFF_972(CK,g1809,g29438);
  dff DFF_973(CK,g1807,g29439);
  dff DFF_974(CK,g1810,g27700);
  dff DFF_975(CK,g1813,g27701);
  dff DFF_976(CK,g1816,g27702);
  dff DFF_977(CK,g1819,g27703);
  dff DFF_978(CK,g1822,g27704);
  dff DFF_979(CK,g1825,g27705);
  dff DFF_980(CK,g1829,g28684);
  dff DFF_981(CK,g1830,g28685);
  dff DFF_982(CK,g1828,g28686);
  dff DFF_983(CK,g1693,g29803);
  dff DFF_984(CK,g1694,g29804);
  dff DFF_985(CK,g1695,g29805);
  dff DFF_986(CK,g1696,g30887);
  dff DFF_987(CK,g1697,g30888);
  dff DFF_988(CK,g1698,g30889);
  dff DFF_989(CK,g1699,g30716);
  dff DFF_990(CK,g1700,g30717);
  dff DFF_991(CK,g1701,g30718);
  dff DFF_992(CK,g1703,g29642);
  dff DFF_993(CK,g1704,g29643);
  dff DFF_994(CK,g1702,g29644);
  dff DFF_995(CK,g1784,g27221);
  dff DFF_996(CK,g1785,g27222);
  dff DFF_997(CK,g1783,g27223);
  dff DFF_998(CK,g1831,g11563);
  dff DFF_999(CK,g1832,g1831);
  dff DFF_1000(CK,g1833,g11564);
  dff DFF_1001(CK,g1834,g1833);
  dff DFF_1002(CK,g1835,g11565);
  dff DFF_1003(CK,g1660,g1835);
  dff DFF_1004(CK,g1661,g11545);
  dff DFF_1005(CK,g1662,g1661);
  dff DFF_1006(CK,g1663,g11546);
  dff DFF_1007(CK,g1664,g1663);
  dff DFF_1008(CK,g1665,g11547);
  dff DFF_1009(CK,g1666,g1665);
  dff DFF_1010(CK,g1667,g11548);
  dff DFF_1011(CK,g1668,g1667);
  dff DFF_1012(CK,g1669,g11549);
  dff DFF_1013(CK,g1670,g1669);
  dff DFF_1014(CK,g1671,g13439);
  dff DFF_1015(CK,g1672,g1671);
  dff DFF_1016(CK,g1680,g19036);
  dff DFF_1017(CK,g1686,g29428);
  dff DFF_1018(CK,g1689,g29429);
  dff DFF_1019(CK,g1678,g29430);
  dff DFF_1020(CK,g1677,g29431);
  dff DFF_1021(CK,g1676,g29432);
  dff DFF_1022(CK,g1675,g29433);
  dff DFF_1023(CK,g1685,g19040);
  dff DFF_1024(CK,g1684,g19039);
  dff DFF_1025(CK,g1683,g19038);
  dff DFF_1026(CK,g1682,g19037);
  dff DFF_1027(CK,g1681,g25152);
  dff DFF_1028(CK,g1679,g27220);
  dff DFF_1029(CK,g1723,g11551);
  dff DFF_1030(CK,g1730,g1723);
  dff DFF_1031(CK,g1731,g11552);
  dff DFF_1032(CK,g1732,g1731);
  dff DFF_1033(CK,g1733,g11553);
  dff DFF_1034(CK,g1734,g1733);
  dff DFF_1035(CK,g1738,g11554);
  dff DFF_1036(CK,g1745,g1738);
  dff DFF_1037(CK,g1746,g11555);
  dff DFF_1038(CK,g1747,g1746);
  dff DFF_1039(CK,g1748,g11556);
  dff DFF_1040(CK,g1749,g1748);
  dff DFF_1041(CK,g1753,g11557);
  dff DFF_1042(CK,g1760,g1753);
  dff DFF_1043(CK,g1761,g11558);
  dff DFF_1044(CK,g1762,g1761);
  dff DFF_1045(CK,g1763,g11559);
  dff DFF_1046(CK,g1764,g1763);
  dff DFF_1047(CK,g1768,g11560);
  dff DFF_1048(CK,g1775,g1768);
  dff DFF_1049(CK,g1776,g11561);
  dff DFF_1050(CK,g1777,g1776);
  dff DFF_1051(CK,g1778,g11562);
  dff DFF_1052(CK,g1705,g1778);
  dff DFF_1053(CK,g1706,g13440);
  dff DFF_1054(CK,g1712,g1706);
  dff DFF_1055(CK,g1718,g1712);
  dff DFF_1056(CK,g1925,g13451);
  dff DFF_1057(CK,g1931,g1925);
  dff DFF_1058(CK,g1930,g1931);
  dff DFF_1059(CK,g1934,g23236);
  dff DFF_1060(CK,g1937,g20564);
  dff DFF_1061(CK,g1890,g20565);
  dff DFF_1062(CK,g1893,g16471);
  dff DFF_1063(CK,g1903,g1893);
  dff DFF_1064(CK,g1904,g1903);
  dff DFF_1065(CK,g1944,g11566);
  dff DFF_1066(CK,g1949,g1944);
  dff DFF_1067(CK,g1950,g11569);
  dff DFF_1068(CK,g1951,g1950);
  dff DFF_1069(CK,g1952,g11570);
  dff DFF_1070(CK,g1953,g1952);
  dff DFF_1071(CK,g1954,g11571);
  dff DFF_1072(CK,g1945,g1954);
  dff DFF_1073(CK,g1946,g11567);
  dff DFF_1074(CK,g1947,g1946);
  dff DFF_1075(CK,g1948,g11568);
  dff DFF_1076(CK,g1870,g1948);
  dff DFF_1077(CK,g1855,g13441);
  dff DFF_1078(CK,g1862,g1855);
  dff DFF_1079(CK,g1866,g1862);
  dff DFF_1080(CK,g1867,g24374);
  dff DFF_1081(CK,g1868,g24375);
  dff DFF_1082(CK,g1869,g24376);
  dff DFF_1083(CK,g1836,g25161);
  dff DFF_1084(CK,g1839,g25153);
  dff DFF_1085(CK,g1842,g25154);
  dff DFF_1086(CK,g1858,g25158);
  dff DFF_1087(CK,g1859,g25159);
  dff DFF_1088(CK,g1860,g25160);
  dff DFF_1089(CK,g1861,g24371);
  dff DFF_1090(CK,g1865,g24372);
  dff DFF_1091(CK,g1845,g24373);
  dff DFF_1092(CK,g1846,g25155);
  dff DFF_1093(CK,g1849,g25156);
  dff DFF_1094(CK,g1852,g25157);
  dff DFF_1095(CK,g1908,g16472);
  dff DFF_1096(CK,g1915,g1908);
  dff DFF_1097(CK,g1922,g1915);
  dff DFF_1098(CK,g1923,g19045);
  dff DFF_1099(CK,g1924,g1923);
  dff DFF_1100(CK,g1928,g29445);
  dff DFF_1101(CK,g1929,g19046);
  dff DFF_1102(CK,g1880,g1929);
  dff DFF_1103(CK,g1938,g19047);
  dff DFF_1104(CK,g1939,g1938);
  dff DFF_1105(CK,g1956,g28271);
  dff DFF_1106(CK,g1957,g28272);
  dff DFF_1107(CK,g1955,g28273);
  dff DFF_1108(CK,g1959,g28274);
  dff DFF_1109(CK,g1960,g28275);
  dff DFF_1110(CK,g1958,g28276);
  dff DFF_1111(CK,g1962,g28277);
  dff DFF_1112(CK,g1963,g28278);
  dff DFF_1113(CK,g1961,g28279);
  dff DFF_1114(CK,g1965,g28280);
  dff DFF_1115(CK,g1966,g28281);
  dff DFF_1116(CK,g1964,g28282);
  dff DFF_1117(CK,g1967,g26003);
  dff DFF_1118(CK,g1970,g26004);
  dff DFF_1119(CK,g1973,g26005);
  dff DFF_1120(CK,g1976,g26006);
  dff DFF_1121(CK,g1979,g26007);
  dff DFF_1122(CK,g1982,g26008);
  dff DFF_1123(CK,g1994,g29151);
  dff DFF_1124(CK,g1997,g29152);
  dff DFF_1125(CK,g2000,g29153);
  dff DFF_1126(CK,g1985,g29148);
  dff DFF_1127(CK,g1988,g29149);
  dff DFF_1128(CK,g1991,g29150);
  dff DFF_1129(CK,g1871,g27224);
  dff DFF_1130(CK,g1874,g27225);
  dff DFF_1131(CK,g1877,g27226);
  dff DFF_1132(CK,g1886,g8302);
  dff DFF_1133(CK,g1887,g24377);
  dff DFF_1134(CK,g1888,g19041);
  dff DFF_1135(CK,g1889,g19042);
  dff DFF_1136(CK,g1894,g19043);
  dff DFF_1137(CK,g1895,g19044);
  dff DFF_1138(CK,g1896,g29444);
  dff DFF_1139(CK,g1897,g29443);
  dff DFF_1140(CK,g1898,g29442);
  dff DFF_1141(CK,g1899,g29441);
  dff DFF_1142(CK,g1900,g29440);
  dff DFF_1143(CK,g1905,g1900);
  dff DFF_1144(CK,g1909,g13442);
  dff DFF_1145(CK,g1910,g13443);
  dff DFF_1146(CK,g1911,g13444);
  dff DFF_1147(CK,g1912,g13445);
  dff DFF_1148(CK,g1913,g13446);
  dff DFF_1149(CK,g1914,g13447);
  dff DFF_1150(CK,g1916,g13448);
  dff DFF_1151(CK,g1917,g13449);
  dff DFF_1152(CK,g1918,g26002);
  dff DFF_1153(CK,g1921,g13450);
  dff DFF_1154(CK,g2003,g13452);
  dff DFF_1155(CK,g2006,g2003);
  dff DFF_1156(CK,g2009,g2006);
  dff DFF_1157(CK,g2010,g20566);
  dff DFF_1158(CK,g2039,g21945);
  dff DFF_1159(CK,g2020,g23237);
  dff DFF_1160(CK,g2013,g24378);
  dff DFF_1161(CK,g2033,g25162);
  dff DFF_1162(CK,g2026,g26009);
  dff DFF_1163(CK,g2040,g26725);
  dff DFF_1164(CK,g2052,g27227);
  dff DFF_1165(CK,g2046,g27706);
  dff DFF_1166(CK,g2059,g28283);
  dff DFF_1167(CK,g2066,g28687);
  dff DFF_1168(CK,g2072,g29154);
  dff DFF_1169(CK,g2079,g23238);
  dff DFF_1170(CK,g2080,g23239);
  dff DFF_1171(CK,g2078,g23240);
  dff DFF_1172(CK,g2082,g23241);
  dff DFF_1173(CK,g2083,g23242);
  dff DFF_1174(CK,g2081,g23243);
  dff DFF_1175(CK,g2085,g23244);
  dff DFF_1176(CK,g2086,g23245);
  dff DFF_1177(CK,g2084,g23246);
  dff DFF_1178(CK,g2088,g23247);
  dff DFF_1179(CK,g2089,g23248);
  dff DFF_1180(CK,g2087,g23249);
  dff DFF_1181(CK,g2091,g23250);
  dff DFF_1182(CK,g2092,g23251);
  dff DFF_1183(CK,g2090,g23252);
  dff DFF_1184(CK,g2094,g23253);
  dff DFF_1185(CK,g2095,g23254);
  dff DFF_1186(CK,g2093,g23255);
  dff DFF_1187(CK,g2097,g23256);
  dff DFF_1188(CK,g2098,g23257);
  dff DFF_1189(CK,g2096,g23258);
  dff DFF_1190(CK,g2100,g23259);
  dff DFF_1191(CK,g2101,g23260);
  dff DFF_1192(CK,g2099,g23261);
  dff DFF_1193(CK,g2103,g23262);
  dff DFF_1194(CK,g2104,g23263);
  dff DFF_1195(CK,g2102,g23264);
  dff DFF_1196(CK,g2106,g23265);
  dff DFF_1197(CK,g2107,g23266);
  dff DFF_1198(CK,g2105,g23267);
  dff DFF_1199(CK,g2109,g23268);
  dff DFF_1200(CK,g2110,g23269);
  dff DFF_1201(CK,g2108,g23270);
  dff DFF_1202(CK,g2112,g23271);
  dff DFF_1203(CK,g2113,g23272);
  dff DFF_1204(CK,g2111,g23273);
  dff DFF_1205(CK,g2115,g26726);
  dff DFF_1206(CK,g2116,g26727);
  dff DFF_1207(CK,g2114,g26728);
  dff DFF_1208(CK,g2118,g24379);
  dff DFF_1209(CK,g2119,g24380);
  dff DFF_1210(CK,g2117,g24381);
  dff DFF_1211(CK,g2214,g13453);
  dff DFF_1212(CK,g2211,g2214);
  dff DFF_1213(CK,g2241,g2211);
  dff DFF_1214(CK,g2206,g24382);
  dff DFF_1215(CK,g2207,g24383);
  dff DFF_1216(CK,g2205,g24384);
  dff DFF_1217(CK,g2209,g24385);
  dff DFF_1218(CK,g2210,g24386);
  dff DFF_1219(CK,g2208,g24387);
  dff DFF_1220(CK,g2218,g24388);
  dff DFF_1221(CK,g2219,g24389);
  dff DFF_1222(CK,g2217,g24390);
  dff DFF_1223(CK,g2221,g24391);
  dff DFF_1224(CK,g2222,g24392);
  dff DFF_1225(CK,g2220,g24393);
  dff DFF_1226(CK,g2224,g24394);
  dff DFF_1227(CK,g2225,g24395);
  dff DFF_1228(CK,g2223,g24396);
  dff DFF_1229(CK,g2227,g24397);
  dff DFF_1230(CK,g2228,g24398);
  dff DFF_1231(CK,g2226,g24399);
  dff DFF_1232(CK,g2230,g24400);
  dff DFF_1233(CK,g2231,g24401);
  dff DFF_1234(CK,g2229,g24402);
  dff DFF_1235(CK,g2233,g24403);
  dff DFF_1236(CK,g2234,g24404);
  dff DFF_1237(CK,g2232,g24405);
  dff DFF_1238(CK,g2236,g24406);
  dff DFF_1239(CK,g2237,g24407);
  dff DFF_1240(CK,g2235,g24408);
  dff DFF_1241(CK,g2239,g24409);
  dff DFF_1242(CK,g2240,g24410);
  dff DFF_1243(CK,g2238,g24411);
  dff DFF_1244(CK,g2245,g26730);
  dff DFF_1245(CK,g2246,g26731);
  dff DFF_1246(CK,g2244,g26732);
  dff DFF_1247(CK,g2248,g26733);
  dff DFF_1248(CK,g2249,g26734);
  dff DFF_1249(CK,g2247,g26735);
  dff DFF_1250(CK,g2251,g26736);
  dff DFF_1251(CK,g2252,g26737);
  dff DFF_1252(CK,g2250,g26738);
  dff DFF_1253(CK,g2254,g26739);
  dff DFF_1254(CK,g2255,g26740);
  dff DFF_1255(CK,g2253,g26741);
  dff DFF_1256(CK,g2261,g30551);
  dff DFF_1257(CK,g2264,g30552);
  dff DFF_1258(CK,g2267,g30553);
  dff DFF_1259(CK,g2306,g30896);
  dff DFF_1260(CK,g2309,g30897);
  dff DFF_1261(CK,g2312,g30898);
  dff DFF_1262(CK,g2270,g30890);
  dff DFF_1263(CK,g2273,g30891);
  dff DFF_1264(CK,g2276,g30892);
  dff DFF_1265(CK,g2315,g30899);
  dff DFF_1266(CK,g2318,g30900);
  dff DFF_1267(CK,g2321,g30901);
  dff DFF_1268(CK,g2279,g30554);
  dff DFF_1269(CK,g2282,g30555);
  dff DFF_1270(CK,g2285,g30556);
  dff DFF_1271(CK,g2324,g30560);
  dff DFF_1272(CK,g2327,g30561);
  dff DFF_1273(CK,g2330,g30562);
  dff DFF_1274(CK,g2288,g30557);
  dff DFF_1275(CK,g2291,g30558);
  dff DFF_1276(CK,g2294,g30559);
  dff DFF_1277(CK,g2333,g30563);
  dff DFF_1278(CK,g2336,g30564);
  dff DFF_1279(CK,g2339,g30565);
  dff DFF_1280(CK,g2297,g30893);
  dff DFF_1281(CK,g2300,g30894);
  dff DFF_1282(CK,g2303,g30895);
  dff DFF_1283(CK,g2342,g30902);
  dff DFF_1284(CK,g2345,g30903);
  dff DFF_1285(CK,g2348,g30904);
  dff DFF_1286(CK,g2160,g26010);
  dff DFF_1287(CK,g2156,g26729);
  dff DFF_1288(CK,g2151,g27228);
  dff DFF_1289(CK,g2147,g27707);
  dff DFF_1290(CK,g2142,g28284);
  dff DFF_1291(CK,g2138,g28688);
  dff DFF_1292(CK,g2133,g29155);
  dff DFF_1293(CK,g2129,g29446);
  dff DFF_1294(CK,g2124,g29648);
  dff DFF_1295(CK,g2120,g29806);
  dff DFF_1296(CK,g2256,g20567);
  dff DFF_1297(CK,g2258,g2256);
  dff DFF_1298(CK,g2257,g2258);
  dff DFF_1299(CK,g2351,g13454);
  dff DFF_1300(CK,g2480,g2351);
  dff DFF_1301(CK,g2476,g2480);
  dff DFF_1302(CK,g2384,g11577);
  dff DFF_1303(CK,g2429,g28285);
  dff DFF_1304(CK,g2418,g28286);
  dff DFF_1305(CK,g2421,g28287);
  dff DFF_1306(CK,g2444,g28288);
  dff DFF_1307(CK,g2433,g28289);
  dff DFF_1308(CK,g2436,g28290);
  dff DFF_1309(CK,g2459,g28291);
  dff DFF_1310(CK,g2448,g28292);
  dff DFF_1311(CK,g2451,g28293);
  dff DFF_1312(CK,g2473,g28294);
  dff DFF_1313(CK,g2463,g28295);
  dff DFF_1314(CK,g2466,g28296);
  dff DFF_1315(CK,g2483,g29447);
  dff DFF_1316(CK,g2486,g29448);
  dff DFF_1317(CK,g2489,g29449);
  dff DFF_1318(CK,g2492,g29652);
  dff DFF_1319(CK,g2495,g29653);
  dff DFF_1320(CK,g2498,g29654);
  dff DFF_1321(CK,g2502,g29450);
  dff DFF_1322(CK,g2503,g29451);
  dff DFF_1323(CK,g2501,g29452);
  dff DFF_1324(CK,g2504,g27708);
  dff DFF_1325(CK,g2507,g27709);
  dff DFF_1326(CK,g2510,g27710);
  dff DFF_1327(CK,g2513,g27711);
  dff DFF_1328(CK,g2516,g27712);
  dff DFF_1329(CK,g2519,g27713);
  dff DFF_1330(CK,g2523,g28689);
  dff DFF_1331(CK,g2524,g28690);
  dff DFF_1332(CK,g2522,g28691);
  dff DFF_1333(CK,g2387,g29807);
  dff DFF_1334(CK,g2388,g29808);
  dff DFF_1335(CK,g2389,g29809);
  dff DFF_1336(CK,g2390,g30905);
  dff DFF_1337(CK,g2391,g30906);
  dff DFF_1338(CK,g2392,g30907);
  dff DFF_1339(CK,g2393,g30719);
  dff DFF_1340(CK,g2394,g30720);
  dff DFF_1341(CK,g2395,g30721);
  dff DFF_1342(CK,g2397,g29649);
  dff DFF_1343(CK,g2398,g29650);
  dff DFF_1344(CK,g2396,g29651);
  dff DFF_1345(CK,g2478,g27230);
  dff DFF_1346(CK,g2479,g27231);
  dff DFF_1347(CK,g2477,g27232);
  dff DFF_1348(CK,g2525,g11590);
  dff DFF_1349(CK,g2526,g2525);
  dff DFF_1350(CK,g2527,g11591);
  dff DFF_1351(CK,g2528,g2527);
  dff DFF_1352(CK,g2529,g11592);
  dff DFF_1353(CK,g2354,g2529);
  dff DFF_1354(CK,g2355,g11572);
  dff DFF_1355(CK,g2356,g2355);
  dff DFF_1356(CK,g2357,g11573);
  dff DFF_1357(CK,g2358,g2357);
  dff DFF_1358(CK,g2359,g11574);
  dff DFF_1359(CK,g2360,g2359);
  dff DFF_1360(CK,g2361,g11575);
  dff DFF_1361(CK,g2362,g2361);
  dff DFF_1362(CK,g2363,g11576);
  dff DFF_1363(CK,g2364,g2363);
  dff DFF_1364(CK,g2365,g13455);
  dff DFF_1365(CK,g2366,g2365);
  dff DFF_1366(CK,g2374,g19048);
  dff DFF_1367(CK,g2380,g30314);
  dff DFF_1368(CK,g2383,g30315);
  dff DFF_1369(CK,g2372,g30316);
  dff DFF_1370(CK,g2371,g30317);
  dff DFF_1371(CK,g2370,g30318);
  dff DFF_1372(CK,g2369,g30319);
  dff DFF_1373(CK,g2379,g19052);
  dff DFF_1374(CK,g2378,g19051);
  dff DFF_1375(CK,g2377,g19050);
  dff DFF_1376(CK,g2376,g19049);
  dff DFF_1377(CK,g2375,g25163);
  dff DFF_1378(CK,g2373,g27229);
  dff DFF_1379(CK,g2417,g11578);
  dff DFF_1380(CK,g2424,g2417);
  dff DFF_1381(CK,g2425,g11579);
  dff DFF_1382(CK,g2426,g2425);
  dff DFF_1383(CK,g2427,g11580);
  dff DFF_1384(CK,g2428,g2427);
  dff DFF_1385(CK,g2432,g11581);
  dff DFF_1386(CK,g2439,g2432);
  dff DFF_1387(CK,g2440,g11582);
  dff DFF_1388(CK,g2441,g2440);
  dff DFF_1389(CK,g2442,g11583);
  dff DFF_1390(CK,g2443,g2442);
  dff DFF_1391(CK,g2447,g11584);
  dff DFF_1392(CK,g2454,g2447);
  dff DFF_1393(CK,g2455,g11585);
  dff DFF_1394(CK,g2456,g2455);
  dff DFF_1395(CK,g2457,g11586);
  dff DFF_1396(CK,g2458,g2457);
  dff DFF_1397(CK,g2462,g11587);
  dff DFF_1398(CK,g2469,g2462);
  dff DFF_1399(CK,g2470,g11588);
  dff DFF_1400(CK,g2471,g2470);
  dff DFF_1401(CK,g2472,g11589);
  dff DFF_1402(CK,g2399,g2472);
  dff DFF_1403(CK,g2400,g13456);
  dff DFF_1404(CK,g2406,g2400);
  dff DFF_1405(CK,g2412,g2406);
  dff DFF_1406(CK,g2619,g13467);
  dff DFF_1407(CK,g2625,g2619);
  dff DFF_1408(CK,g2624,g2625);
  dff DFF_1409(CK,g2628,g23274);
  dff DFF_1410(CK,g2631,g20568);
  dff DFF_1411(CK,g2584,g20569);
  dff DFF_1412(CK,g2587,g16473);
  dff DFF_1413(CK,g2597,g2587);
  dff DFF_1414(CK,g2598,g2597);
  dff DFF_1415(CK,g2638,g11593);
  dff DFF_1416(CK,g2643,g2638);
  dff DFF_1417(CK,g2644,g11596);
  dff DFF_1418(CK,g2645,g2644);
  dff DFF_1419(CK,g2646,g11597);
  dff DFF_1420(CK,g2647,g2646);
  dff DFF_1421(CK,g2648,g11598);
  dff DFF_1422(CK,g2639,g2648);
  dff DFF_1423(CK,g2640,g11594);
  dff DFF_1424(CK,g2641,g2640);
  dff DFF_1425(CK,g2642,g11595);
  dff DFF_1426(CK,g2564,g2642);
  dff DFF_1427(CK,g2549,g13457);
  dff DFF_1428(CK,g2556,g2549);
  dff DFF_1429(CK,g2560,g2556);
  dff DFF_1430(CK,g2561,g24415);
  dff DFF_1431(CK,g2562,g24416);
  dff DFF_1432(CK,g2563,g24417);
  dff DFF_1433(CK,g2530,g25172);
  dff DFF_1434(CK,g2533,g25164);
  dff DFF_1435(CK,g2536,g25165);
  dff DFF_1436(CK,g2552,g25169);
  dff DFF_1437(CK,g2553,g25170);
  dff DFF_1438(CK,g2554,g25171);
  dff DFF_1439(CK,g2555,g24412);
  dff DFF_1440(CK,g2559,g24413);
  dff DFF_1441(CK,g2539,g24414);
  dff DFF_1442(CK,g2540,g25166);
  dff DFF_1443(CK,g2543,g25167);
  dff DFF_1444(CK,g2546,g25168);
  dff DFF_1445(CK,g2602,g16474);
  dff DFF_1446(CK,g2609,g2602);
  dff DFF_1447(CK,g2616,g2609);
  dff DFF_1448(CK,g2617,g19057);
  dff DFF_1449(CK,g2618,g2617);
  dff DFF_1450(CK,g2622,g30325);
  dff DFF_1451(CK,g2623,g19058);
  dff DFF_1452(CK,g2574,g2623);
  dff DFF_1453(CK,g2632,g19059);
  dff DFF_1454(CK,g2633,g2632);
  dff DFF_1455(CK,g2650,g28297);
  dff DFF_1456(CK,g2651,g28298);
  dff DFF_1457(CK,g2649,g28299);
  dff DFF_1458(CK,g2653,g28300);
  dff DFF_1459(CK,g2654,g28301);
  dff DFF_1460(CK,g2652,g28302);
  dff DFF_1461(CK,g2656,g28303);
  dff DFF_1462(CK,g2657,g28304);
  dff DFF_1463(CK,g2655,g28305);
  dff DFF_1464(CK,g2659,g28306);
  dff DFF_1465(CK,g2660,g28307);
  dff DFF_1466(CK,g2658,g28308);
  dff DFF_1467(CK,g2661,g26012);
  dff DFF_1468(CK,g2664,g26013);
  dff DFF_1469(CK,g2667,g26014);
  dff DFF_1470(CK,g2670,g26015);
  dff DFF_1471(CK,g2673,g26016);
  dff DFF_1472(CK,g2676,g26017);
  dff DFF_1473(CK,g2688,g29159);
  dff DFF_1474(CK,g2691,g29160);
  dff DFF_1475(CK,g2694,g29161);
  dff DFF_1476(CK,g2679,g29156);
  dff DFF_1477(CK,g2682,g29157);
  dff DFF_1478(CK,g2685,g29158);
  dff DFF_1479(CK,g2565,g27233);
  dff DFF_1480(CK,g2568,g27234);
  dff DFF_1481(CK,g2571,g27235);
  dff DFF_1482(CK,g2580,g8311);
  dff DFF_1483(CK,g2581,g24418);
  dff DFF_1484(CK,g2582,g19053);
  dff DFF_1485(CK,g2583,g19054);
  dff DFF_1486(CK,g2588,g19055);
  dff DFF_1487(CK,g2589,g19056);
  dff DFF_1488(CK,g2590,g30324);
  dff DFF_1489(CK,g2591,g30323);
  dff DFF_1490(CK,g2592,g30322);
  dff DFF_1491(CK,g2593,g30321);
  dff DFF_1492(CK,g2594,g30320);
  dff DFF_1493(CK,g2599,g2594);
  dff DFF_1494(CK,g2603,g13458);
  dff DFF_1495(CK,g2604,g13459);
  dff DFF_1496(CK,g2605,g13460);
  dff DFF_1497(CK,g2606,g13461);
  dff DFF_1498(CK,g2607,g13462);
  dff DFF_1499(CK,g2608,g13463);
  dff DFF_1500(CK,g2610,g13464);
  dff DFF_1501(CK,g2611,g13465);
  dff DFF_1502(CK,g2612,g26011);
  dff DFF_1503(CK,g2615,g13466);
  dff DFF_1504(CK,g2697,g13468);
  dff DFF_1505(CK,g2700,g2697);
  dff DFF_1506(CK,g2703,g2700);
  dff DFF_1507(CK,g2704,g20570);
  dff DFF_1508(CK,g2733,g21946);
  dff DFF_1509(CK,g2714,g23275);
  dff DFF_1510(CK,g2707,g24419);
  dff DFF_1511(CK,g2727,g25173);
  dff DFF_1512(CK,g2720,g26018);
  dff DFF_1513(CK,g2734,g26742);
  dff DFF_1514(CK,g2746,g27236);
  dff DFF_1515(CK,g2740,g27714);
  dff DFF_1516(CK,g2753,g28309);
  dff DFF_1517(CK,g2760,g28692);
  dff DFF_1518(CK,g2766,g29162);
  dff DFF_1519(CK,g2773,g23276);
  dff DFF_1520(CK,g2774,g23277);
  dff DFF_1521(CK,g2772,g23278);
  dff DFF_1522(CK,g2776,g23279);
  dff DFF_1523(CK,g2777,g23280);
  dff DFF_1524(CK,g2775,g23281);
  dff DFF_1525(CK,g2779,g23282);
  dff DFF_1526(CK,g2780,g23283);
  dff DFF_1527(CK,g2778,g23284);
  dff DFF_1528(CK,g2782,g23285);
  dff DFF_1529(CK,g2783,g23286);
  dff DFF_1530(CK,g2781,g23287);
  dff DFF_1531(CK,g2785,g23288);
  dff DFF_1532(CK,g2786,g23289);
  dff DFF_1533(CK,g2784,g23290);
  dff DFF_1534(CK,g2788,g23291);
  dff DFF_1535(CK,g2789,g23292);
  dff DFF_1536(CK,g2787,g23293);
  dff DFF_1537(CK,g2791,g23294);
  dff DFF_1538(CK,g2792,g23295);
  dff DFF_1539(CK,g2790,g23296);
  dff DFF_1540(CK,g2794,g23297);
  dff DFF_1541(CK,g2795,g23298);
  dff DFF_1542(CK,g2793,g23299);
  dff DFF_1543(CK,g2797,g23300);
  dff DFF_1544(CK,g2798,g23301);
  dff DFF_1545(CK,g2796,g23302);
  dff DFF_1546(CK,g2800,g23303);
  dff DFF_1547(CK,g2801,g23304);
  dff DFF_1548(CK,g2799,g23305);
  dff DFF_1549(CK,g2803,g23306);
  dff DFF_1550(CK,g2804,g23307);
  dff DFF_1551(CK,g2802,g23308);
  dff DFF_1552(CK,g2806,g23309);
  dff DFF_1553(CK,g2807,g23310);
  dff DFF_1554(CK,g2805,g23311);
  dff DFF_1555(CK,g2809,g26743);
  dff DFF_1556(CK,g2810,g26744);
  dff DFF_1557(CK,g2808,g26745);
  dff DFF_1558(CK,g2812,g24420);
  dff DFF_1559(CK,g2813,g24421);
  dff DFF_1560(CK,g2811,g24422);
  dff DFF_1561(CK,g3054,g23317);
  dff DFF_1562(CK,g3079,g23318);
  dff DFF_1563(CK,g3080,g21965);
  dff DFF_1564(CK,g3043,g29453);
  dff DFF_1565(CK,g3044,g29454);
  dff DFF_1566(CK,g3045,g29455);
  dff DFF_1567(CK,g3046,g29456);
  dff DFF_1568(CK,g3047,g29457);
  dff DFF_1569(CK,g3048,g29458);
  dff DFF_1570(CK,g3049,g29459);
  dff DFF_1571(CK,g3050,g29460);
  dff DFF_1572(CK,g3051,g29655);
  dff DFF_1573(CK,g3052,g29972);
  dff DFF_1574(CK,g3053,g29973);
  dff DFF_1575(CK,g3055,g29974);
  dff DFF_1576(CK,g3056,g29975);
  dff DFF_1577(CK,g3057,g29976);
  dff DFF_1578(CK,g3058,g29977);
  dff DFF_1579(CK,g3059,g29978);
  dff DFF_1580(CK,g3060,g29979);
  dff DFF_1581(CK,g3061,g30119);
  dff DFF_1582(CK,g3062,g30908);
  dff DFF_1583(CK,g3063,g30909);
  dff DFF_1584(CK,g3064,g30910);
  dff DFF_1585(CK,g3065,g30911);
  dff DFF_1586(CK,g3066,g30912);
  dff DFF_1587(CK,g3067,g30913);
  dff DFF_1588(CK,g3068,g30914);
  dff DFF_1589(CK,g3069,g30915);
  dff DFF_1590(CK,g3070,g30940);
  dff DFF_1591(CK,g3071,g30980);
  dff DFF_1592(CK,g3072,g30981);
  dff DFF_1593(CK,g3073,g30982);
  dff DFF_1594(CK,g3074,g30983);
  dff DFF_1595(CK,g3075,g30984);
  dff DFF_1596(CK,g3076,g30985);
  dff DFF_1597(CK,g3077,g30986);
  dff DFF_1598(CK,g3078,g30987);
  dff DFF_1599(CK,g2997,g30989);
  dff DFF_1600(CK,g2993,g26748);
  dff DFF_1601(CK,g2998,g27238);
  dff DFF_1602(CK,g3006,g25177);
  dff DFF_1603(CK,g3002,g26021);
  dff DFF_1604(CK,g3013,g26750);
  dff DFF_1605(CK,g3010,g27239);
  dff DFF_1606(CK,g3024,g27716);
  dff DFF_1607(CK,g3018,g24425);
  dff DFF_1608(CK,g3028,g25176);
  dff DFF_1609(CK,g3036,g26022);
  dff DFF_1610(CK,g3032,g26749);
  dff DFF_1611(CK,g3040,g16497);
  dff DFF_1612(CK,g2986,g3040);
  dff DFF_1613(CK,g2987,g16495);
  dff DFF_1614(CK,g48,g20595);
  dff DFF_1615(CK,g45,g20596);
  dff DFF_1616(CK,g42,g20597);
  dff DFF_1617(CK,g39,g20598);
  dff DFF_1618(CK,g27,g20599);
  dff DFF_1619(CK,g30,g20600);
  dff DFF_1620(CK,g33,g20601);
  dff DFF_1621(CK,g36,g20602);
  dff DFF_1622(CK,g3083,g20603);
  dff DFF_1623(CK,g26,g20604);
  dff DFF_1624(CK,g2992,g21966);
  dff DFF_1625(CK,g23,g20605);
  dff DFF_1626(CK,g20,g20606);
  dff DFF_1627(CK,g17,g20607);
  dff DFF_1628(CK,g11,g20608);
  dff DFF_1629(CK,g14,g20589);
  dff DFF_1630(CK,g5,g20590);
  dff DFF_1631(CK,g8,g20591);
  dff DFF_1632(CK,g2,g20592);
  dff DFF_1633(CK,g2990,g20593);
  dff DFF_1634(CK,g2991,g21964);
  dff DFF_1635(CK,g1,g20594);
  not NOT_0(II13089,g563);
  not NOT_1(g562,II13089);
  not NOT_2(II13092,g1249);
  not NOT_3(g1248,II13092);
  not NOT_4(II13095,g1943);
  not NOT_5(g1942,II13095);
  not NOT_6(II13098,g2637);
  not NOT_7(g2636,II13098);
  not NOT_8(II13101,g1);
  not NOT_9(g3235,II13101);
  not NOT_10(II13104,g2);
  not NOT_11(g3236,II13104);
  not NOT_12(II13107,g5);
  not NOT_13(g3237,II13107);
  not NOT_14(II13110,g8);
  not NOT_15(g3238,II13110);
  not NOT_16(II13113,g11);
  not NOT_17(g3239,II13113);
  not NOT_18(II13116,g14);
  not NOT_19(g3240,II13116);
  not NOT_20(II13119,g17);
  not NOT_21(g3241,II13119);
  not NOT_22(II13122,g20);
  not NOT_23(g3242,II13122);
  not NOT_24(II13125,g23);
  not NOT_25(g3243,II13125);
  not NOT_26(II13128,g26);
  not NOT_27(g3244,II13128);
  not NOT_28(II13131,g27);
  not NOT_29(g3245,II13131);
  not NOT_30(II13134,g30);
  not NOT_31(g3246,II13134);
  not NOT_32(II13137,g33);
  not NOT_33(g3247,II13137);
  not NOT_34(II13140,g36);
  not NOT_35(g3248,II13140);
  not NOT_36(II13143,g39);
  not NOT_37(g3249,II13143);
  not NOT_38(II13146,g42);
  not NOT_39(g3250,II13146);
  not NOT_40(II13149,g45);
  not NOT_41(g3251,II13149);
  not NOT_42(II13152,g48);
  not NOT_43(g3252,II13152);
  not NOT_44(II13155,g51);
  not NOT_45(g3253,II13155);
  not NOT_46(II13158,g165);
  not NOT_47(g3254,II13158);
  not NOT_48(II13161,g308);
  not NOT_49(g3304,II13161);
  not NOT_50(g3305,g305);
  not NOT_51(II13165,g401);
  not NOT_52(g3306,II13165);
  not NOT_53(g3337,g309);
  not NOT_54(II13169,g550);
  not NOT_55(g3338,II13169);
  not NOT_56(g3365,g499);
  not NOT_57(II13173,g629);
  not NOT_58(g3366,II13173);
  not NOT_59(II13176,g630);
  not NOT_60(g3398,II13176);
  not NOT_61(II13179,g853);
  not NOT_62(g3410,II13179);
  not NOT_63(II13182,g995);
  not NOT_64(g3460,II13182);
  not NOT_65(g3461,g992);
  not NOT_66(II13186,g1088);
  not NOT_67(g3462,II13186);
  not NOT_68(g3493,g996);
  not NOT_69(II13190,g1236);
  not NOT_70(g3494,II13190);
  not NOT_71(g3521,g1186);
  not NOT_72(II13194,g1315);
  not NOT_73(g3522,II13194);
  not NOT_74(II13197,g1316);
  not NOT_75(g3554,II13197);
  not NOT_76(II13200,g1547);
  not NOT_77(g3566,II13200);
  not NOT_78(II13203,g1689);
  not NOT_79(g3616,II13203);
  not NOT_80(g3617,g1686);
  not NOT_81(II13207,g1782);
  not NOT_82(g3618,II13207);
  not NOT_83(g3649,g1690);
  not NOT_84(II13211,g1930);
  not NOT_85(g3650,II13211);
  not NOT_86(g3677,g1880);
  not NOT_87(II13215,g2009);
  not NOT_88(g3678,II13215);
  not NOT_89(II13218,g2010);
  not NOT_90(g3710,II13218);
  not NOT_91(II13221,g2241);
  not NOT_92(g3722,II13221);
  not NOT_93(II13224,g2383);
  not NOT_94(g3772,II13224);
  not NOT_95(g3773,g2380);
  not NOT_96(II13228,g2476);
  not NOT_97(g3774,II13228);
  not NOT_98(g3805,g2384);
  not NOT_99(II13232,g2624);
  not NOT_100(g3806,II13232);
  not NOT_101(g3833,g2574);
  not NOT_102(II13236,g2703);
  not NOT_103(g3834,II13236);
  not NOT_104(II13239,g2704);
  not NOT_105(g3866,II13239);
  not NOT_106(II13242,g2879);
  not NOT_107(g3878,II13242);
  not NOT_108(g3897,g2950);
  not NOT_109(II13246,g2987);
  not NOT_110(g3900,II13246);
  not NOT_111(g3919,g3080);
  not NOT_112(g3922,g150);
  not NOT_113(g3925,g155);
  not NOT_114(g3928,g157);
  not NOT_115(g3931,g171);
  not NOT_116(g3934,g176);
  not NOT_117(g3937,g178);
  not NOT_118(g3940,g408);
  not NOT_119(g3941,g455);
  not NOT_120(g3942,g699);
  not NOT_121(g3945,g726);
  not NOT_122(g3948,g835);
  not NOT_123(g3951,g840);
  not NOT_124(g3954,g842);
  not NOT_125(g3957,g856);
  not NOT_126(g3960,g861);
  not NOT_127(g3963,g863);
  not NOT_128(g3966,g1526);
  not NOT_129(g3969,g1531);
  not NOT_130(g3972,g1533);
  not NOT_131(g3975,g1552);
  not NOT_132(g3978,g1554);
  not NOT_133(g3981,g2217);
  not NOT_134(g3984,g2222);
  not NOT_135(g3987,g2224);
  not NOT_136(g3990,g2245);
  not NOT_137(II13275,g2848);
  not NOT_138(g3993,II13275);
  not NOT_139(g3994,g2848);
  not NOT_140(g3995,g3064);
  not NOT_141(g3996,g3073);
  not NOT_142(g3997,g45);
  not NOT_143(g3998,g23);
  not NOT_144(g3999,g3204);
  not NOT_145(g4000,g153);
  not NOT_146(g4003,g158);
  not NOT_147(g4006,g160);
  not NOT_148(g4009,g174);
  not NOT_149(g4012,g179);
  not NOT_150(g4015,g411);
  not NOT_151(g4016,g417);
  not NOT_152(g4017,g427);
  not NOT_153(g4020,g700);
  not NOT_154(g4023,g702);
  not NOT_155(g4026,g727);
  not NOT_156(g4029,g838);
  not NOT_157(g4032,g843);
  not NOT_158(g4035,g845);
  not NOT_159(g4038,g859);
  not NOT_160(g4041,g864);
  not NOT_161(g4044,g866);
  not NOT_162(g4047,g1095);
  not NOT_163(g4048,g1142);
  not NOT_164(g4049,g1385);
  not NOT_165(g4052,g1412);
  not NOT_166(g4055,g1529);
  not NOT_167(g4058,g1534);
  not NOT_168(g4061,g1536);
  not NOT_169(g4064,g1550);
  not NOT_170(g4067,g1555);
  not NOT_171(g4070,g1557);
  not NOT_172(g4073,g2220);
  not NOT_173(g4076,g2225);
  not NOT_174(g4079,g2227);
  not NOT_175(g4082,g2246);
  not NOT_176(g4085,g2248);
  not NOT_177(II13316,g2836);
  not NOT_178(g4088,II13316);
  not NOT_179(g4089,g2836);
  not NOT_180(II13320,g2864);
  not NOT_181(g4090,II13320);
  not NOT_182(g4091,g2864);
  not NOT_183(g4092,g3074);
  not NOT_184(g4093,g33);
  not NOT_185(g4094,g3207);
  not NOT_186(g4095,g130);
  not NOT_187(g4098,g156);
  not NOT_188(g4101,g161);
  not NOT_189(g4104,g163);
  not NOT_190(g4107,g177);
  not NOT_191(g4110,g414);
  not NOT_192(g4111,g420);
  not NOT_193(g4112,g428);
  not NOT_194(g4115,g698);
  not NOT_195(g4118,g703);
  not NOT_196(g4121,g705);
  not NOT_197(g4124,g725);
  not NOT_198(g4127,g841);
  not NOT_199(g4130,g846);
  not NOT_200(g4133,g848);
  not NOT_201(g4136,g862);
  not NOT_202(g4139,g867);
  not NOT_203(g4142,g1098);
  not NOT_204(g4143,g1104);
  not NOT_205(g4144,g1114);
  not NOT_206(g4147,g1386);
  not NOT_207(g4150,g1388);
  not NOT_208(g4153,g1413);
  not NOT_209(g4156,g1532);
  not NOT_210(g4159,g1537);
  not NOT_211(g4162,g1539);
  not NOT_212(g4165,g1553);
  not NOT_213(g4168,g1558);
  not NOT_214(g4171,g1560);
  not NOT_215(g4174,g1789);
  not NOT_216(g4175,g1836);
  not NOT_217(g4176,g2079);
  not NOT_218(g4179,g2106);
  not NOT_219(g4182,g2223);
  not NOT_220(g4185,g2228);
  not NOT_221(g4188,g2230);
  not NOT_222(g4191,g2244);
  not NOT_223(g4194,g2249);
  not NOT_224(g4197,g2251);
  not NOT_225(II13366,g2851);
  not NOT_226(g4200,II13366);
  not NOT_227(g4201,g2851);
  not NOT_228(g4202,g42);
  not NOT_229(g4203,g20);
  not NOT_230(g4204,g3188);
  not NOT_231(g4205,g131);
  not NOT_232(g4208,g133);
  not NOT_233(g4211,g159);
  not NOT_234(g4214,g164);
  not NOT_235(g4217,g354);
  not NOT_236(g4220,g423);
  not NOT_237(g4221,g426);
  not NOT_238(g4224,g429);
  not NOT_239(g4225,g701);
  not NOT_240(g4228,g706);
  not NOT_241(g4231,g708);
  not NOT_242(g4234,g818);
  not NOT_243(g4237,g844);
  not NOT_244(g4240,g849);
  not NOT_245(g4243,g851);
  not NOT_246(g4246,g865);
  not NOT_247(g4249,g1101);
  not NOT_248(g4250,g1107);
  not NOT_249(g4251,g1115);
  not NOT_250(g4254,g1384);
  not NOT_251(g4257,g1389);
  not NOT_252(g4260,g1391);
  not NOT_253(g4263,g1411);
  not NOT_254(g4266,g1535);
  not NOT_255(g4269,g1540);
  not NOT_256(g4272,g1542);
  not NOT_257(g4275,g1556);
  not NOT_258(g4278,g1561);
  not NOT_259(g4281,g1792);
  not NOT_260(g4282,g1798);
  not NOT_261(g4283,g1808);
  not NOT_262(g4286,g2080);
  not NOT_263(g4289,g2082);
  not NOT_264(g4292,g2107);
  not NOT_265(g4295,g2226);
  not NOT_266(g4298,g2231);
  not NOT_267(g4301,g2233);
  not NOT_268(g4304,g2247);
  not NOT_269(g4307,g2252);
  not NOT_270(g4310,g2254);
  not NOT_271(g4313,g2483);
  not NOT_272(g4314,g2530);
  not NOT_273(g4315,g2773);
  not NOT_274(g4318,g2800);
  not NOT_275(II13417,g2839);
  not NOT_276(g4321,II13417);
  not NOT_277(g4322,g2839);
  not NOT_278(II13421,g2867);
  not NOT_279(g4323,II13421);
  not NOT_280(g4324,g2867);
  not NOT_281(g4325,g36);
  not NOT_282(g4326,g181);
  not NOT_283(g4329,g129);
  not NOT_284(g4332,g134);
  not NOT_285(g4335,g162);
  not NOT_286(II13430,g101);
  not NOT_287(g4338,II13430);
  not NOT_288(II13433,g105);
  not NOT_289(g4339,II13433);
  not NOT_290(g4340,g343);
  not NOT_291(g4343,g369);
  not NOT_292(g4346,g432);
  not NOT_293(g4347,g438);
  not NOT_294(g4348,g704);
  not NOT_295(g4351,g709);
  not NOT_296(g4354,g711);
  not NOT_297(g4357,g729);
  not NOT_298(g4360,g819);
  not NOT_299(g4363,g821);
  not NOT_300(g4366,g847);
  not NOT_301(g4369,g852);
  not NOT_302(g4372,g1041);
  not NOT_303(g4375,g1110);
  not NOT_304(g4376,g1113);
  not NOT_305(g4379,g1116);
  not NOT_306(g4380,g1387);
  not NOT_307(g4383,g1392);
  not NOT_308(g4386,g1394);
  not NOT_309(g4389,g1512);
  not NOT_310(g4392,g1538);
  not NOT_311(g4395,g1543);
  not NOT_312(g4398,g1545);
  not NOT_313(g4401,g1559);
  not NOT_314(g4404,g1795);
  not NOT_315(g4405,g1801);
  not NOT_316(g4406,g1809);
  not NOT_317(g4409,g2078);
  not NOT_318(g4412,g2083);
  not NOT_319(g4415,g2085);
  not NOT_320(g4418,g2105);
  not NOT_321(g4421,g2229);
  not NOT_322(g4424,g2234);
  not NOT_323(g4427,g2236);
  not NOT_324(g4430,g2250);
  not NOT_325(g4433,g2255);
  not NOT_326(g4436,g2486);
  not NOT_327(g4437,g2492);
  not NOT_328(g4438,g2502);
  not NOT_329(g4441,g2774);
  not NOT_330(g4444,g2776);
  not NOT_331(g4447,g2801);
  not NOT_332(II13478,g2854);
  not NOT_333(g4450,II13478);
  not NOT_334(g4451,g2854);
  not NOT_335(g4452,g17);
  not NOT_336(g4453,g132);
  not NOT_337(g4456,g309);
  not NOT_338(g4465,g346);
  not NOT_339(g4468,g358);
  not NOT_340(g4471,g384);
  not NOT_341(g4474,g435);
  not NOT_342(g4475,g441);
  not NOT_343(g4476,g576);
  not NOT_344(g4479,g587);
  not NOT_345(g4480,g707);
  not NOT_346(g4483,g712);
  not NOT_347(g4486,g714);
  not NOT_348(g4489,g730);
  not NOT_349(g4492,g732);
  not NOT_350(g4495,g869);
  not NOT_351(g4498,g817);
  not NOT_352(g4501,g822);
  not NOT_353(g4504,g850);
  not NOT_354(II13501,g789);
  not NOT_355(g4507,II13501);
  not NOT_356(II13504,g793);
  not NOT_357(g4508,II13504);
  not NOT_358(g4509,g1030);
  not NOT_359(g4512,g1056);
  not NOT_360(g4515,g1119);
  not NOT_361(g4516,g1125);
  not NOT_362(g4517,g1390);
  not NOT_363(g4520,g1395);
  not NOT_364(g4523,g1397);
  not NOT_365(g4526,g1415);
  not NOT_366(g4529,g1513);
  not NOT_367(g4532,g1515);
  not NOT_368(g4535,g1541);
  not NOT_369(g4538,g1546);
  not NOT_370(g4541,g1735);
  not NOT_371(g4544,g1804);
  not NOT_372(g4545,g1807);
  not NOT_373(g4548,g1810);
  not NOT_374(g4549,g2081);
  not NOT_375(g4552,g2086);
  not NOT_376(g4555,g2088);
  not NOT_377(g4558,g2206);
  not NOT_378(g4561,g2232);
  not NOT_379(g4564,g2237);
  not NOT_380(g4567,g2239);
  not NOT_381(g4570,g2253);
  not NOT_382(g4573,g2489);
  not NOT_383(g4574,g2495);
  not NOT_384(g4575,g2503);
  not NOT_385(g4578,g2772);
  not NOT_386(g4581,g2777);
  not NOT_387(g4584,g2779);
  not NOT_388(g4587,g2799);
  not NOT_389(II13538,g2870);
  not NOT_390(g4590,II13538);
  not NOT_391(g4591,g2870);
  not NOT_392(g4592,g361);
  not NOT_393(g4595,g373);
  not NOT_394(g4598,g398);
  not NOT_395(g4601,g444);
  not NOT_396(g4602,g525);
  not NOT_397(g4603,g577);
  not NOT_398(g4606,g579);
  not NOT_399(g4609,g590);
  not NOT_400(g4610,g596);
  not NOT_401(g4611,g710);
  not NOT_402(g4614,g715);
  not NOT_403(g4617,g717);
  not NOT_404(g4620,g728);
  not NOT_405(g4623,g733);
  not NOT_406(g4626,g735);
  not NOT_407(g4629,g820);
  not NOT_408(g4632,g996);
  not NOT_409(g4641,g1033);
  not NOT_410(g4644,g1045);
  not NOT_411(g4647,g1071);
  not NOT_412(g4650,g1122);
  not NOT_413(g4651,g1128);
  not NOT_414(g4652,g1262);
  not NOT_415(g4655,g1273);
  not NOT_416(g4656,g1393);
  not NOT_417(g4659,g1398);
  not NOT_418(g4662,g1400);
  not NOT_419(g4665,g1416);
  not NOT_420(g4668,g1418);
  not NOT_421(g4671,g1563);
  not NOT_422(g4674,g1511);
  not NOT_423(g4677,g1516);
  not NOT_424(g4680,g1544);
  not NOT_425(II13575,g1476);
  not NOT_426(g4683,II13575);
  not NOT_427(II13578,g1481);
  not NOT_428(g4684,II13578);
  not NOT_429(g4685,g1724);
  not NOT_430(g4688,g1750);
  not NOT_431(g4691,g1813);
  not NOT_432(g4692,g1819);
  not NOT_433(g4693,g2084);
  not NOT_434(g4696,g2089);
  not NOT_435(g4699,g2091);
  not NOT_436(g4702,g2109);
  not NOT_437(g4705,g2207);
  not NOT_438(g4708,g2209);
  not NOT_439(g4711,g2235);
  not NOT_440(g4714,g2240);
  not NOT_441(g4717,g2429);
  not NOT_442(g4720,g2498);
  not NOT_443(g4721,g2501);
  not NOT_444(g4724,g2504);
  not NOT_445(g4725,g2775);
  not NOT_446(g4728,g2780);
  not NOT_447(g4731,g2782);
  not NOT_448(g4734,g11);
  not NOT_449(II13601,g121);
  not NOT_450(g4735,II13601);
  not NOT_451(II13604,g125);
  not NOT_452(g4736,II13604);
  not NOT_453(g4737,g376);
  not NOT_454(g4740,g388);
  not NOT_455(g4743,g575);
  not NOT_456(g4746,g580);
  not NOT_457(g4749,g582);
  not NOT_458(g4752,g593);
  not NOT_459(g4753,g599);
  not NOT_460(g4754,g713);
  not NOT_461(g4757,g718);
  not NOT_462(g4760,g720);
  not NOT_463(g4763,g731);
  not NOT_464(g4766,g736);
  not NOT_465(g4769,g1048);
  not NOT_466(g4772,g1060);
  not NOT_467(g4775,g1085);
  not NOT_468(g4778,g1131);
  not NOT_469(g4779,g1211);
  not NOT_470(g4780,g1263);
  not NOT_471(g4783,g1265);
  not NOT_472(g4786,g1276);
  not NOT_473(g4787,g1282);
  not NOT_474(g4788,g1396);
  not NOT_475(g4791,g1401);
  not NOT_476(g4794,g1403);
  not NOT_477(g4797,g1414);
  not NOT_478(g4800,g1419);
  not NOT_479(g4803,g1421);
  not NOT_480(g4806,g1514);
  not NOT_481(g4809,g1690);
  not NOT_482(g4818,g1727);
  not NOT_483(g4821,g1739);
  not NOT_484(g4824,g1765);
  not NOT_485(g4827,g1816);
  not NOT_486(g4828,g1822);
  not NOT_487(g4829,g1956);
  not NOT_488(g4832,g1967);
  not NOT_489(g4833,g2087);
  not NOT_490(g4836,g2092);
  not NOT_491(g4839,g2094);
  not NOT_492(g4842,g2110);
  not NOT_493(g4845,g2112);
  not NOT_494(g4848,g2257);
  not NOT_495(g4851,g2205);
  not NOT_496(g4854,g2210);
  not NOT_497(g4857,g2238);
  not NOT_498(II13652,g2170);
  not NOT_499(g4860,II13652);
  not NOT_500(II13655,g2175);
  not NOT_501(g4861,II13655);
  not NOT_502(g4862,g2418);
  not NOT_503(g4865,g2444);
  not NOT_504(g4868,g2507);
  not NOT_505(g4869,g2513);
  not NOT_506(g4870,g2778);
  not NOT_507(g4873,g2783);
  not NOT_508(g4876,g2785);
  not NOT_509(g4879,g2803);
  not NOT_510(g4882,g391);
  not NOT_511(g4885,g448);
  not NOT_512(g4888,g578);
  not NOT_513(g4891,g583);
  not NOT_514(g4894,g585);
  not NOT_515(g4897,g602);
  not NOT_516(g4898,g605);
  not NOT_517(g4899,g716);
  not NOT_518(g4902,g721);
  not NOT_519(g4905,g723);
  not NOT_520(g4908,g734);
  not NOT_521(II13677,g809);
  not NOT_522(g4911,II13677);
  not NOT_523(II13680,g813);
  not NOT_524(g4912,II13680);
  not NOT_525(g4913,g1063);
  not NOT_526(g4916,g1075);
  not NOT_527(g4919,g1261);
  not NOT_528(g4922,g1266);
  not NOT_529(g4925,g1268);
  not NOT_530(g4928,g1279);
  not NOT_531(g4929,g1285);
  not NOT_532(g4930,g1399);
  not NOT_533(g4933,g1404);
  not NOT_534(g4936,g1406);
  not NOT_535(g4939,g1417);
  not NOT_536(g4942,g1422);
  not NOT_537(g4945,g1742);
  not NOT_538(g4948,g1754);
  not NOT_539(g4951,g1779);
  not NOT_540(g4954,g1825);
  not NOT_541(g4955,g1905);
  not NOT_542(g4956,g1957);
  not NOT_543(g4959,g1959);
  not NOT_544(g4962,g1970);
  not NOT_545(g4963,g1976);
  not NOT_546(g4964,g2090);
  not NOT_547(g4967,g2095);
  not NOT_548(g4970,g2097);
  not NOT_549(g4973,g2108);
  not NOT_550(g4976,g2113);
  not NOT_551(g4979,g2115);
  not NOT_552(g4982,g2208);
  not NOT_553(g4985,g2384);
  not NOT_554(g4994,g2421);
  not NOT_555(g4997,g2433);
  not NOT_556(g5000,g2459);
  not NOT_557(g5003,g2510);
  not NOT_558(g5004,g2516);
  not NOT_559(g5005,g2650);
  not NOT_560(g5008,g2661);
  not NOT_561(g5009,g2781);
  not NOT_562(g5012,g2786);
  not NOT_563(g5015,g2788);
  not NOT_564(g5018,g2804);
  not NOT_565(g5021,g2806);
  not NOT_566(g5024,g449);
  not NOT_567(g5027,g581);
  not NOT_568(g5030,g586);
  not NOT_569(g5033,g608);
  not NOT_570(g5034,g614);
  not NOT_571(g5035,g719);
  not NOT_572(g5038,g724);
  not NOT_573(g5041,g1078);
  not NOT_574(g5044,g1135);
  not NOT_575(g5047,g1264);
  not NOT_576(g5050,g1269);
  not NOT_577(g5053,g1271);
  not NOT_578(g5056,g1288);
  not NOT_579(g5057,g1291);
  not NOT_580(g5058,g1402);
  not NOT_581(g5061,g1407);
  not NOT_582(g5064,g1409);
  not NOT_583(g5067,g1420);
  not NOT_584(II13742,g1501);
  not NOT_585(g5070,II13742);
  not NOT_586(II13745,g1506);
  not NOT_587(g5071,II13745);
  not NOT_588(g5072,g1757);
  not NOT_589(g5075,g1769);
  not NOT_590(g5078,g1955);
  not NOT_591(g5081,g1960);
  not NOT_592(g5084,g1962);
  not NOT_593(g5087,g1973);
  not NOT_594(g5088,g1979);
  not NOT_595(g5089,g2093);
  not NOT_596(g5092,g2098);
  not NOT_597(g5095,g2100);
  not NOT_598(g5098,g2111);
  not NOT_599(g5101,g2116);
  not NOT_600(g5104,g2436);
  not NOT_601(g5107,g2448);
  not NOT_602(g5110,g2473);
  not NOT_603(g5113,g2519);
  not NOT_604(g5114,g2599);
  not NOT_605(g5115,g2651);
  not NOT_606(g5118,g2653);
  not NOT_607(g5121,g2664);
  not NOT_608(g5122,g2670);
  not NOT_609(g5123,g2784);
  not NOT_610(g5126,g2789);
  not NOT_611(g5129,g2791);
  not NOT_612(g5132,g2802);
  not NOT_613(g5135,g2807);
  not NOT_614(g5138,g2809);
  not NOT_615(II13775,g109);
  not NOT_616(g5141,II13775);
  not NOT_617(g5142,g447);
  not NOT_618(g5145,g584);
  not NOT_619(g5148,g611);
  not NOT_620(g5149,g617);
  not NOT_621(g5150,g722);
  not NOT_622(g5153,g1136);
  not NOT_623(g5156,g1267);
  not NOT_624(g5159,g1272);
  not NOT_625(g5162,g1294);
  not NOT_626(g5163,g1300);
  not NOT_627(g5164,g1405);
  not NOT_628(g5167,g1410);
  not NOT_629(g5170,g1772);
  not NOT_630(g5173,g1829);
  not NOT_631(g5176,g1958);
  not NOT_632(g5179,g1963);
  not NOT_633(g5182,g1965);
  not NOT_634(g5185,g1982);
  not NOT_635(g5186,g1985);
  not NOT_636(g5187,g2096);
  not NOT_637(g5190,g2101);
  not NOT_638(g5193,g2103);
  not NOT_639(g5196,g2114);
  not NOT_640(II13801,g2195);
  not NOT_641(g5199,II13801);
  not NOT_642(II13804,g2200);
  not NOT_643(g5200,II13804);
  not NOT_644(g5201,g2451);
  not NOT_645(g5204,g2463);
  not NOT_646(g5207,g2649);
  not NOT_647(g5210,g2654);
  not NOT_648(g5213,g2656);
  not NOT_649(g5216,g2667);
  not NOT_650(g5217,g2673);
  not NOT_651(g5218,g2787);
  not NOT_652(g5221,g2792);
  not NOT_653(g5224,g2794);
  not NOT_654(g5227,g2805);
  not NOT_655(g5230,g2810);
  not NOT_656(g5233,g620);
  not NOT_657(II13820,g797);
  not NOT_658(g5234,II13820);
  not NOT_659(g5235,g1134);
  not NOT_660(g5238,g1270);
  not NOT_661(g5241,g1297);
  not NOT_662(g5242,g1303);
  not NOT_663(g5243,g1408);
  not NOT_664(g5246,g1830);
  not NOT_665(g5249,g1961);
  not NOT_666(g5252,g1966);
  not NOT_667(g5255,g1988);
  not NOT_668(g5256,g1994);
  not NOT_669(g5257,g2099);
  not NOT_670(g5260,g2104);
  not NOT_671(g5263,g2466);
  not NOT_672(g5266,g2523);
  not NOT_673(g5269,g2652);
  not NOT_674(g5272,g2657);
  not NOT_675(g5275,g2659);
  not NOT_676(g5278,g2676);
  not NOT_677(g5279,g2679);
  not NOT_678(g5280,g2790);
  not NOT_679(g5283,g2795);
  not NOT_680(g5286,g2797);
  not NOT_681(g5289,g2808);
  not NOT_682(g5292,g2857);
  not NOT_683(g5293,g738);
  not NOT_684(g5296,g1306);
  not NOT_685(II13849,g1486);
  not NOT_686(g5297,II13849);
  not NOT_687(g5298,g1828);
  not NOT_688(g5301,g1964);
  not NOT_689(g5304,g1991);
  not NOT_690(g5305,g1997);
  not NOT_691(g5306,g2102);
  not NOT_692(g5309,g2524);
  not NOT_693(g5312,g2655);
  not NOT_694(g5315,g2660);
  not NOT_695(g5318,g2682);
  not NOT_696(g5319,g2688);
  not NOT_697(g5320,g2793);
  not NOT_698(g5323,g2798);
  not NOT_699(g5326,g2873);
  not NOT_700(g5327,g739);
  not NOT_701(g5330,g1424);
  not NOT_702(g5333,g2000);
  not NOT_703(II13868,g2180);
  not NOT_704(g5334,II13868);
  not NOT_705(g5335,g2522);
  not NOT_706(g5338,g2658);
  not NOT_707(g5341,g2685);
  not NOT_708(g5342,g2691);
  not NOT_709(g5343,g2796);
  not NOT_710(g5346,g3106);
  not NOT_711(g5349,g2877);
  not NOT_712(g5352,g737);
  not NOT_713(g5355,g1425);
  not NOT_714(g5358,g2118);
  not NOT_715(g5361,g2694);
  not NOT_716(g5362,g2817);
  not NOT_717(g5363,g3107);
  not NOT_718(g5366,g2878);
  not NOT_719(g5369,g1423);
  not NOT_720(g5372,g2119);
  not NOT_721(g5375,g2812);
  not NOT_722(g5378,g2933);
  not NOT_723(g5379,g3108);
  not NOT_724(g5382,g2117);
  not NOT_725(g5385,g2813);
  not NOT_726(II13892,g3040);
  not NOT_727(g5388,II13892);
  not NOT_728(g5389,g3040);
  not NOT_729(II13896,g343);
  not NOT_730(g5390,II13896);
  not NOT_731(g5391,g2811);
  not NOT_732(g5394,g3054);
  not NOT_733(II13901,g346);
  not NOT_734(g5395,II13901);
  not NOT_735(II13904,g358);
  not NOT_736(g5396,II13904);
  not NOT_737(II13907,g1030);
  not NOT_738(g5397,II13907);
  not NOT_739(II13910,g361);
  not NOT_740(g5398,II13910);
  not NOT_741(II13913,g373);
  not NOT_742(g5399,II13913);
  not NOT_743(II13916,g1033);
  not NOT_744(g5400,II13916);
  not NOT_745(II13919,g1045);
  not NOT_746(g5401,II13919);
  not NOT_747(II13922,g1724);
  not NOT_748(g5402,II13922);
  not NOT_749(II13925,g376);
  not NOT_750(g5403,II13925);
  not NOT_751(II13928,g388);
  not NOT_752(g5404,II13928);
  not NOT_753(II13931,g1048);
  not NOT_754(g5405,II13931);
  not NOT_755(II13934,g1060);
  not NOT_756(g5406,II13934);
  not NOT_757(II13937,g1727);
  not NOT_758(g5407,II13937);
  not NOT_759(II13940,g1739);
  not NOT_760(g5408,II13940);
  not NOT_761(II13943,g2418);
  not NOT_762(g5409,II13943);
  not NOT_763(g5410,g3079);
  not NOT_764(II13947,g391);
  not NOT_765(g5411,II13947);
  not NOT_766(II13950,g1063);
  not NOT_767(g5412,II13950);
  not NOT_768(II13953,g1075);
  not NOT_769(g5413,II13953);
  not NOT_770(II13956,g1742);
  not NOT_771(g5414,II13956);
  not NOT_772(II13959,g1754);
  not NOT_773(g5415,II13959);
  not NOT_774(II13962,g2421);
  not NOT_775(g5416,II13962);
  not NOT_776(II13965,g2433);
  not NOT_777(g5417,II13965);
  not NOT_778(II13968,g1078);
  not NOT_779(g5418,II13968);
  not NOT_780(II13971,g1757);
  not NOT_781(g5419,II13971);
  not NOT_782(II13974,g1769);
  not NOT_783(g5420,II13974);
  not NOT_784(II13977,g2436);
  not NOT_785(g5421,II13977);
  not NOT_786(II13980,g2448);
  not NOT_787(g5422,II13980);
  not NOT_788(g5423,g2879);
  not NOT_789(II13984,g1772);
  not NOT_790(g5424,II13984);
  not NOT_791(II13987,g2451);
  not NOT_792(g5425,II13987);
  not NOT_793(II13990,g2463);
  not NOT_794(g5426,II13990);
  not NOT_795(II13993,g2466);
  not NOT_796(g5427,II13993);
  not NOT_797(g5428,g3210);
  not NOT_798(g5431,g3211);
  not NOT_799(g5434,g3084);
  not NOT_800(II13999,g276);
  not NOT_801(g5437,II13999);
  not NOT_802(II14002,g276);
  not NOT_803(g5438,II14002);
  not NOT_804(g5469,g3085);
  not NOT_805(II14006,g963);
  not NOT_806(g5472,II14006);
  not NOT_807(II14009,g963);
  not NOT_808(g5473,II14009);
  not NOT_809(g5504,g3086);
  not NOT_810(g5507,g3155);
  not NOT_811(II14014,g499);
  not NOT_812(g5508,II14014);
  not NOT_813(II14017,g1657);
  not NOT_814(g5511,II14017);
  not NOT_815(II14020,g1657);
  not NOT_816(g5512,II14020);
  not NOT_817(g5543,g3087);
  not NOT_818(g5546,g3164);
  not NOT_819(g5547,g101);
  not NOT_820(g5548,g105);
  not NOT_821(II14027,g182);
  not NOT_822(g5549,II14027);
  not NOT_823(II14030,g182);
  not NOT_824(g5550,II14030);
  not NOT_825(g5551,g514);
  not NOT_826(II14034,g1186);
  not NOT_827(g5552,II14034);
  not NOT_828(II14037,g2351);
  not NOT_829(g5555,II14037);
  not NOT_830(II14040,g2351);
  not NOT_831(g5556,II14040);
  not NOT_832(g5587,g3091);
  not NOT_833(g5590,g3158);
  not NOT_834(g5591,g3173);
  not NOT_835(g5592,g515);
  not NOT_836(g5593,g789);
  not NOT_837(g5594,g793);
  not NOT_838(II14049,g870);
  not NOT_839(g5595,II14049);
  not NOT_840(II14052,g870);
  not NOT_841(g5596,II14052);
  not NOT_842(g5597,g1200);
  not NOT_843(II14056,g1880);
  not NOT_844(g5598,II14056);
  not NOT_845(g5601,g3092);
  not NOT_846(g5604,g3167);
  not NOT_847(g5605,g3182);
  not NOT_848(g5606,g79);
  not NOT_849(g5609,g1201);
  not NOT_850(g5610,g1476);
  not NOT_851(g5611,g1481);
  not NOT_852(II14066,g1564);
  not NOT_853(g5612,II14066);
  not NOT_854(II14069,g1564);
  not NOT_855(g5613,II14069);
  not NOT_856(g5614,g1894);
  not NOT_857(II14073,g2574);
  not NOT_858(g5615,II14073);
  not NOT_859(g5618,g3093);
  not NOT_860(g5621,g3161);
  not NOT_861(g5622,g3176);
  not NOT_862(g5623,g70);
  not NOT_863(g5626,g121);
  not NOT_864(g5627,g125);
  not NOT_865(g5628,g300);
  not NOT_866(II14083,g325);
  not NOT_867(g5629,II14083);
  not NOT_868(g5631,g767);
  not NOT_869(g5634,g1895);
  not NOT_870(g5635,g2170);
  not NOT_871(g5636,g2175);
  not NOT_872(II14091,g2258);
  not NOT_873(g5637,II14091);
  not NOT_874(II14094,g2258);
  not NOT_875(g5638,II14094);
  not NOT_876(g5639,g2588);
  not NOT_877(g5640,g3170);
  not NOT_878(g5641,g3185);
  not NOT_879(g5642,g61);
  not NOT_880(g5645,g101);
  not NOT_881(g5646,g213);
  not NOT_882(g5647,g301);
  not NOT_883(II14104,g331);
  not NOT_884(g5648,II14104);
  not NOT_885(g5651,g758);
  not NOT_886(g5654,g809);
  not NOT_887(g5655,g813);
  not NOT_888(g5656,g987);
  not NOT_889(II14113,g1012);
  not NOT_890(g5657,II14113);
  not NOT_891(g5659,g1453);
  not NOT_892(g5662,g2589);
  not NOT_893(g5663,g3179);
  not NOT_894(g5664,g65);
  not NOT_895(g5665,g105);
  not NOT_896(g5666,g216);
  not NOT_897(g5667,g222);
  not NOT_898(g5668,g299);
  not NOT_899(g5675,g302);
  not NOT_900(g5679,g506);
  not NOT_901(g5680,g749);
  not NOT_902(g5683,g789);
  not NOT_903(g5684,g900);
  not NOT_904(g5685,g988);
  not NOT_905(II14134,g1018);
  not NOT_906(g5686,II14134);
  not NOT_907(g5689,g1444);
  not NOT_908(g5692,g1501);
  not NOT_909(g5693,g1506);
  not NOT_910(g5694,g1681);
  not NOT_911(II14143,g1706);
  not NOT_912(g5695,II14143);
  not NOT_913(g5697,g2147);
  not NOT_914(g5700,g3088);
  not NOT_915(II14149,g3231);
  not NOT_916(g5701,II14149);
  not NOT_917(g5702,g56);
  not NOT_918(g5703,g109);
  not NOT_919(g5704,g219);
  not NOT_920(g5705,g225);
  not NOT_921(g5706,g231);
  not NOT_922(g5707,g109);
  not NOT_923(g5708,g303);
  not NOT_924(g5712,g305);
  not NOT_925(II14163,g113);
  not NOT_926(g5713,II14163);
  not NOT_927(g5714,g507);
  not NOT_928(g5715,g541);
  not NOT_929(g5716,g753);
  not NOT_930(g5717,g793);
  not NOT_931(g5718,g903);
  not NOT_932(g5719,g909);
  not NOT_933(g5720,g986);
  not NOT_934(g5727,g989);
  not NOT_935(g5731,g1192);
  not NOT_936(g5732,g1435);
  not NOT_937(g5735,g1476);
  not NOT_938(g5736,g1594);
  not NOT_939(g5737,g1682);
  not NOT_940(II14182,g1712);
  not NOT_941(g5738,II14182);
  not NOT_942(g5741,g2138);
  not NOT_943(g5744,g2195);
  not NOT_944(g5745,g2200);
  not NOT_945(g5746,g2375);
  not NOT_946(II14191,g2400);
  not NOT_947(g5747,II14191);
  not NOT_948(II14195,g3212);
  not NOT_949(g5749,II14195);
  not NOT_950(g5750,g92);
  not NOT_951(g5751,g52);
  not NOT_952(g5752,g113);
  not NOT_953(g5753,g228);
  not NOT_954(g5754,g234);
  not NOT_955(g5755,g240);
  not NOT_956(g5756,g304);
  not NOT_957(g5759,g508);
  not NOT_958(g5760,g744);
  not NOT_959(g5761,g797);
  not NOT_960(g5762,g906);
  not NOT_961(g5763,g912);
  not NOT_962(g5764,g918);
  not NOT_963(g5765,g797);
  not NOT_964(g5766,g990);
  not NOT_965(g5770,g992);
  not NOT_966(II14219,g801);
  not NOT_967(g5771,II14219);
  not NOT_968(g5772,g1193);
  not NOT_969(g5773,g1227);
  not NOT_970(g5774,g1439);
  not NOT_971(g5775,g1481);
  not NOT_972(g5776,g1597);
  not NOT_973(g5777,g1603);
  not NOT_974(g5778,g1680);
  not NOT_975(g5785,g1683);
  not NOT_976(g5789,g1886);
  not NOT_977(g5790,g2129);
  not NOT_978(g5793,g2170);
  not NOT_979(g5794,g2288);
  not NOT_980(g5795,g2376);
  not NOT_981(II14238,g2406);
  not NOT_982(g5796,II14238);
  not NOT_983(II14243,g3221);
  not NOT_984(g5799,II14243);
  not NOT_985(II14246,g3227);
  not NOT_986(g5800,II14246);
  not NOT_987(II14249,g3216);
  not NOT_988(g5801,II14249);
  not NOT_989(g5802,g83);
  not NOT_990(g5803,g117);
  not NOT_991(g5804,g237);
  not NOT_992(g5805,g243);
  not NOT_993(g5806,g249);
  not NOT_994(g5808,g509);
  not NOT_995(g5809,g780);
  not NOT_996(g5810,g740);
  not NOT_997(g5811,g801);
  not NOT_998(g5812,g915);
  not NOT_999(g5813,g921);
  not NOT_1000(g5814,g927);
  not NOT_1001(g5815,g991);
  not NOT_1002(g5818,g1194);
  not NOT_1003(g5819,g1430);
  not NOT_1004(g5820,g1486);
  not NOT_1005(g5821,g1600);
  not NOT_1006(g5822,g1606);
  not NOT_1007(g5823,g1612);
  not NOT_1008(g5824,g1486);
  not NOT_1009(g5825,g1684);
  not NOT_1010(g5829,g1686);
  not NOT_1011(II14280,g1491);
  not NOT_1012(g5830,II14280);
  not NOT_1013(g5831,g1887);
  not NOT_1014(g5832,g1921);
  not NOT_1015(g5833,g2133);
  not NOT_1016(g5834,g2175);
  not NOT_1017(g5835,g2291);
  not NOT_1018(g5836,g2297);
  not NOT_1019(g5837,g2374);
  not NOT_1020(g5844,g2377);
  not NOT_1021(g5848,g2580);
  not NOT_1022(II14295,g3228);
  not NOT_1023(g5849,II14295);
  not NOT_1024(II14298,g3217);
  not NOT_1025(g5850,II14298);
  not NOT_1026(g5851,g74);
  not NOT_1027(g5852,g121);
  not NOT_1028(g5853,g246);
  not NOT_1029(g5854,g252);
  not NOT_1030(g5855,g258);
  not NOT_1031(II14306,g97);
  not NOT_1032(g5856,II14306);
  not NOT_1033(g5857,g538);
  not NOT_1034(g5858,g771);
  not NOT_1035(g5859,g805);
  not NOT_1036(g5860,g924);
  not NOT_1037(g5861,g930);
  not NOT_1038(g5862,g936);
  not NOT_1039(g5864,g1195);
  not NOT_1040(g5865,g1466);
  not NOT_1041(g5866,g1426);
  not NOT_1042(g5867,g1491);
  not NOT_1043(g5868,g1609);
  not NOT_1044(g5869,g1615);
  not NOT_1045(g5870,g1621);
  not NOT_1046(g5871,g1685);
  not NOT_1047(g5874,g1888);
  not NOT_1048(g5875,g2124);
  not NOT_1049(g5876,g2180);
  not NOT_1050(g5877,g2294);
  not NOT_1051(g5878,g2300);
  not NOT_1052(g5879,g2306);
  not NOT_1053(g5880,g2180);
  not NOT_1054(g5881,g2378);
  not NOT_1055(g5885,g2380);
  not NOT_1056(II14338,g2185);
  not NOT_1057(g5886,II14338);
  not NOT_1058(g5887,g2581);
  not NOT_1059(g5888,g2615);
  not NOT_1060(II14343,g3219);
  not NOT_1061(g5889,II14343);
  not NOT_1062(g5890,g88);
  not NOT_1063(g5893,g125);
  not NOT_1064(g5894,g186);
  not NOT_1065(g5895,g255);
  not NOT_1066(g5896,g261);
  not NOT_1067(g5897,g267);
  not NOT_1068(g5898,g762);
  not NOT_1069(g5899,g809);
  not NOT_1070(g5900,g933);
  not NOT_1071(g5901,g939);
  not NOT_1072(g5902,g945);
  not NOT_1073(II14357,g785);
  not NOT_1074(g5903,II14357);
  not NOT_1075(g5904,g1224);
  not NOT_1076(g5905,g1457);
  not NOT_1077(g5906,g1496);
  not NOT_1078(g5907,g1618);
  not NOT_1079(g5908,g1624);
  not NOT_1080(g5909,g1630);
  not NOT_1081(g5911,g1889);
  not NOT_1082(g5912,g2160);
  not NOT_1083(g5913,g2120);
  not NOT_1084(g5914,g2185);
  not NOT_1085(g5915,g2303);
  not NOT_1086(g5916,g2309);
  not NOT_1087(g5917,g2315);
  not NOT_1088(g5918,g2379);
  not NOT_1089(g5921,g2582);
  not NOT_1090(II14378,g3234);
  not NOT_1091(g5922,II14378);
  not NOT_1092(II14381,g3223);
  not NOT_1093(g5923,II14381);
  not NOT_1094(II14384,g3218);
  not NOT_1095(g5924,II14384);
  not NOT_1096(g5925,g189);
  not NOT_1097(g5926,g195);
  not NOT_1098(g5927,g264);
  not NOT_1099(g5928,g270);
  not NOT_1100(g5929,g776);
  not NOT_1101(g5932,g813);
  not NOT_1102(g5933,g873);
  not NOT_1103(g5934,g942);
  not NOT_1104(g5935,g948);
  not NOT_1105(g5936,g954);
  not NOT_1106(g5937,g1448);
  not NOT_1107(g5938,g1501);
  not NOT_1108(g5939,g1627);
  not NOT_1109(g5940,g1633);
  not NOT_1110(g5941,g1639);
  not NOT_1111(II14402,g1471);
  not NOT_1112(g5942,II14402);
  not NOT_1113(g5943,g1918);
  not NOT_1114(g5944,g2151);
  not NOT_1115(g5945,g2190);
  not NOT_1116(g5946,g2312);
  not NOT_1117(g5947,g2318);
  not NOT_1118(g5948,g2324);
  not NOT_1119(g5950,g2583);
  not NOT_1120(II14413,g3233);
  not NOT_1121(g5951,II14413);
  not NOT_1122(II14416,g3222);
  not NOT_1123(g5952,II14416);
  not NOT_1124(g5953,g97);
  not NOT_1125(g5954,g192);
  not NOT_1126(g5955,g198);
  not NOT_1127(g5956,g204);
  not NOT_1128(g5957,g273);
  not NOT_1129(II14424,g117);
  not NOT_1130(g5958,II14424);
  not NOT_1131(g5959,g876);
  not NOT_1132(g5960,g882);
  not NOT_1133(g5961,g951);
  not NOT_1134(g5962,g957);
  not NOT_1135(g5963,g1462);
  not NOT_1136(g5966,g1506);
  not NOT_1137(g5967,g1567);
  not NOT_1138(g5968,g1636);
  not NOT_1139(g5969,g1642);
  not NOT_1140(g5970,g1648);
  not NOT_1141(g5971,g2142);
  not NOT_1142(g5972,g2195);
  not NOT_1143(g5973,g2321);
  not NOT_1144(g5974,g2327);
  not NOT_1145(g5975,g2333);
  not NOT_1146(II14442,g2165);
  not NOT_1147(g5976,II14442);
  not NOT_1148(g5977,g2612);
  not NOT_1149(II14446,g3230);
  not NOT_1150(g5978,II14446);
  not NOT_1151(II14449,g3224);
  not NOT_1152(g5979,II14449);
  not NOT_1153(g5980,g201);
  not NOT_1154(g5981,g207);
  not NOT_1155(g5982,g785);
  not NOT_1156(g5983,g879);
  not NOT_1157(g5984,g885);
  not NOT_1158(g5985,g891);
  not NOT_1159(g5986,g960);
  not NOT_1160(II14459,g805);
  not NOT_1161(g5987,II14459);
  not NOT_1162(g5988,g1570);
  not NOT_1163(g5989,g1576);
  not NOT_1164(g5990,g1645);
  not NOT_1165(g5991,g1651);
  not NOT_1166(g5992,g2156);
  not NOT_1167(g5995,g2200);
  not NOT_1168(g5996,g2261);
  not NOT_1169(g5997,g2330);
  not NOT_1170(g5998,g2336);
  not NOT_1171(g5999,g2342);
  not NOT_1172(II14472,g3080);
  not NOT_1173(g6000,II14472);
  not NOT_1174(II14475,g3225);
  not NOT_1175(g6014,II14475);
  not NOT_1176(II14478,g3213);
  not NOT_1177(g6015,II14478);
  not NOT_1178(g6016,g210);
  not NOT_1179(g6017,g888);
  not NOT_1180(g6018,g894);
  not NOT_1181(g6019,g1471);
  not NOT_1182(g6020,g1573);
  not NOT_1183(g6021,g1579);
  not NOT_1184(g6022,g1585);
  not NOT_1185(g6023,g1654);
  not NOT_1186(II14489,g1496);
  not NOT_1187(g6024,II14489);
  not NOT_1188(g6025,g2264);
  not NOT_1189(g6026,g2270);
  not NOT_1190(g6027,g2339);
  not NOT_1191(g6028,g2345);
  not NOT_1192(II14496,g3226);
  not NOT_1193(g6029,II14496);
  not NOT_1194(II14499,g3214);
  not NOT_1195(g6030,II14499);
  not NOT_1196(II14502,g471);
  not NOT_1197(g6031,II14502);
  not NOT_1198(g6032,g897);
  not NOT_1199(g6033,g1582);
  not NOT_1200(g6034,g1588);
  not NOT_1201(g6035,g2165);
  not NOT_1202(g6036,g2267);
  not NOT_1203(g6037,g2273);
  not NOT_1204(g6038,g2279);
  not NOT_1205(g6039,g2348);
  not NOT_1206(II14513,g2190);
  not NOT_1207(g6040,II14513);
  not NOT_1208(II14516,g3215);
  not NOT_1209(g6041,II14516);
  not NOT_1210(II14519,g1158);
  not NOT_1211(g6042,II14519);
  not NOT_1212(g6043,g1591);
  not NOT_1213(g6044,g2276);
  not NOT_1214(g6045,g2282);
  not NOT_1215(II14525,g1852);
  not NOT_1216(g6046,II14525);
  not NOT_1217(g6047,g2285);
  not NOT_1218(II14529,g3142);
  not NOT_1219(g6048,II14529);
  not NOT_1220(II14532,g354);
  not NOT_1221(g6051,II14532);
  not NOT_1222(II14535,g2546);
  not NOT_1223(g6052,II14535);
  not NOT_1224(II14538,g369);
  not NOT_1225(g6053,II14538);
  not NOT_1226(II14541,g455);
  not NOT_1227(g6054,II14541);
  not NOT_1228(II14544,g1041);
  not NOT_1229(g6055,II14544);
  not NOT_1230(II14547,g384);
  not NOT_1231(g6056,II14547);
  not NOT_1232(II14550,g458);
  not NOT_1233(g6057,II14550);
  not NOT_1234(II14553,g1056);
  not NOT_1235(g6058,II14553);
  not NOT_1236(II14556,g1142);
  not NOT_1237(g6059,II14556);
  not NOT_1238(II14559,g1735);
  not NOT_1239(g6060,II14559);
  not NOT_1240(II14562,g398);
  not NOT_1241(g6061,II14562);
  not NOT_1242(II14565,g461);
  not NOT_1243(g6062,II14565);
  not NOT_1244(II14568,g1071);
  not NOT_1245(g6063,II14568);
  not NOT_1246(II14571,g1145);
  not NOT_1247(g6064,II14571);
  not NOT_1248(II14574,g1750);
  not NOT_1249(g6065,II14574);
  not NOT_1250(II14577,g1836);
  not NOT_1251(g6066,II14577);
  not NOT_1252(II14580,g2429);
  not NOT_1253(g6067,II14580);
  not NOT_1254(g6068,g499);
  not NOT_1255(II14584,g465);
  not NOT_1256(g6079,II14584);
  not NOT_1257(II14587,g1085);
  not NOT_1258(g6080,II14587);
  not NOT_1259(II14590,g1148);
  not NOT_1260(g6081,II14590);
  not NOT_1261(II14593,g1765);
  not NOT_1262(g6082,II14593);
  not NOT_1263(II14596,g1839);
  not NOT_1264(g6083,II14596);
  not NOT_1265(II14599,g2444);
  not NOT_1266(g6084,II14599);
  not NOT_1267(II14602,g2530);
  not NOT_1268(g6085,II14602);
  not NOT_1269(II14605,g468);
  not NOT_1270(g6086,II14605);
  not NOT_1271(g6087,g1186);
  not NOT_1272(II14609,g1152);
  not NOT_1273(g6098,II14609);
  not NOT_1274(II14612,g1779);
  not NOT_1275(g6099,II14612);
  not NOT_1276(II14615,g1842);
  not NOT_1277(g6100,II14615);
  not NOT_1278(II14618,g2459);
  not NOT_1279(g6101,II14618);
  not NOT_1280(II14621,g2533);
  not NOT_1281(g6102,II14621);
  not NOT_1282(II14624,g1155);
  not NOT_1283(g6103,II14624);
  not NOT_1284(g6104,g1880);
  not NOT_1285(II14628,g1846);
  not NOT_1286(g6115,II14628);
  not NOT_1287(II14631,g2473);
  not NOT_1288(g6116,II14631);
  not NOT_1289(II14634,g2536);
  not NOT_1290(g6117,II14634);
  not NOT_1291(II14637,g1849);
  not NOT_1292(g6118,II14637);
  not NOT_1293(g6119,g2574);
  not NOT_1294(II14641,g2540);
  not NOT_1295(g6130,II14641);
  not NOT_1296(II14644,g3142);
  not NOT_1297(g6131,II14644);
  not NOT_1298(II14647,g2543);
  not NOT_1299(g6134,II14647);
  not NOT_1300(II14650,g525);
  not NOT_1301(g6135,II14650);
  not NOT_1302(g6136,g672);
  not NOT_1303(II14654,g3220);
  not NOT_1304(g6139,II14654);
  not NOT_1305(g6140,g524);
  not NOT_1306(g6141,g554);
  not NOT_1307(g6142,g679);
  not NOT_1308(II14660,g1211);
  not NOT_1309(g6145,II14660);
  not NOT_1310(g6146,g1358);
  not NOT_1311(g6149,g3097);
  not NOT_1312(II14665,g3147);
  not NOT_1313(g6153,II14665);
  not NOT_1314(II14668,g3232);
  not NOT_1315(g6156,II14668);
  not NOT_1316(g6157,g686);
  not NOT_1317(g6161,g1210);
  not NOT_1318(g6162,g1240);
  not NOT_1319(g6163,g1365);
  not NOT_1320(II14675,g1905);
  not NOT_1321(g6166,II14675);
  not NOT_1322(g6167,g2052);
  not NOT_1323(g6170,g3098);
  not NOT_1324(g6173,g557);
  not NOT_1325(g6177,g633);
  not NOT_1326(g6180,g692);
  not NOT_1327(g6183,g291);
  not NOT_1328(g6184,g1372);
  not NOT_1329(g6188,g1904);
  not NOT_1330(g6189,g1934);
  not NOT_1331(g6190,g2059);
  not NOT_1332(II14688,g2599);
  not NOT_1333(g6193,II14688);
  not NOT_1334(g6194,g2746);
  not NOT_1335(g6197,g3099);
  not NOT_1336(g6200,g542);
  not NOT_1337(g6201,g646);
  not NOT_1338(g6204,g289);
  not NOT_1339(g6205,g1243);
  not NOT_1340(g6209,g1319);
  not NOT_1341(g6212,g1378);
  not NOT_1342(g6215,g978);
  not NOT_1343(g6216,g2066);
  not NOT_1344(g6220,g2598);
  not NOT_1345(g6221,g2628);
  not NOT_1346(g6222,g2753);
  not NOT_1347(II14704,g2818);
  not NOT_1348(g6225,II14704);
  not NOT_1349(g6226,g2818);
  not NOT_1350(g6227,g3100);
  not NOT_1351(II14709,g3229);
  not NOT_1352(g6230,II14709);
  not NOT_1353(II14712,g138);
  not NOT_1354(g6231,II14712);
  not NOT_1355(II14715,g138);
  not NOT_1356(g6232,II14715);
  not NOT_1357(g6281,g510);
  not NOT_1358(g6284,g640);
  not NOT_1359(g6288,g287);
  not NOT_1360(g6289,g1228);
  not NOT_1361(g6290,g1332);
  not NOT_1362(g6293,g976);
  not NOT_1363(g6294,g1937);
  not NOT_1364(g6298,g2013);
  not NOT_1365(g6301,g2072);
  not NOT_1366(g6304,g1672);
  not NOT_1367(g6305,g2760);
  not NOT_1368(g6309,g14);
  not NOT_1369(g6310,g3101);
  not NOT_1370(II14731,g135);
  not NOT_1371(g6313,II14731);
  not NOT_1372(II14734,g135);
  not NOT_1373(g6314,II14734);
  not NOT_1374(g6363,g653);
  not NOT_1375(g6367,g285);
  not NOT_1376(II14739,g826);
  not NOT_1377(g6368,II14739);
  not NOT_1378(II14742,g826);
  not NOT_1379(g6369,II14742);
  not NOT_1380(g6418,g1196);
  not NOT_1381(g6421,g1326);
  not NOT_1382(g6425,g974);
  not NOT_1383(g6426,g1922);
  not NOT_1384(g6427,g2026);
  not NOT_1385(g6430,g1670);
  not NOT_1386(g6431,g2631);
  not NOT_1387(g6435,g2707);
  not NOT_1388(g6438,g2766);
  not NOT_1389(g6441,g2366);
  not NOT_1390(II14755,g2821);
  not NOT_1391(g6442,II14755);
  not NOT_1392(g6443,g2821);
  not NOT_1393(g6444,g3102);
  not NOT_1394(II14760,g405);
  not NOT_1395(g6447,II14760);
  not NOT_1396(II14763,g405);
  not NOT_1397(g6448,II14763);
  not NOT_1398(II14766,g545);
  not NOT_1399(g6485,II14766);
  not NOT_1400(II14769,g545);
  not NOT_1401(g6486,II14769);
  not NOT_1402(g6512,g544);
  not NOT_1403(g6513,g660);
  not NOT_1404(g6517,g283);
  not NOT_1405(II14775,g823);
  not NOT_1406(g6518,II14775);
  not NOT_1407(II14778,g823);
  not NOT_1408(g6519,II14778);
  not NOT_1409(g6568,g1339);
  not NOT_1410(g6572,g972);
  not NOT_1411(II14783,g1520);
  not NOT_1412(g6573,II14783);
  not NOT_1413(II14786,g1520);
  not NOT_1414(g6574,II14786);
  not NOT_1415(g6623,g1890);
  not NOT_1416(g6626,g2020);
  not NOT_1417(g6630,g1668);
  not NOT_1418(g6631,g2616);
  not NOT_1419(g6632,g2720);
  not NOT_1420(g6635,g2364);
  not NOT_1421(g6636,g1491);
  not NOT_1422(g6637,g5);
  not NOT_1423(g6638,g3103);
  not NOT_1424(g6641,g113);
  not NOT_1425(II14799,g551);
  not NOT_1426(g6642,II14799);
  not NOT_1427(II14802,g551);
  not NOT_1428(g6643,II14802);
  not NOT_1429(g6672,g464);
  not NOT_1430(g6675,g458);
  not NOT_1431(g6676,g559);
  not NOT_1432(II14808,g623);
  not NOT_1433(g6677,II14808);
  not NOT_1434(II14811,g623);
  not NOT_1435(g6678,II14811);
  not NOT_1436(g6707,g666);
  not NOT_1437(g6711,g281);
  not NOT_1438(II14816,g1092);
  not NOT_1439(g6712,II14816);
  not NOT_1440(II14819,g1092);
  not NOT_1441(g6713,II14819);
  not NOT_1442(II14822,g1231);
  not NOT_1443(g6750,II14822);
  not NOT_1444(II14825,g1231);
  not NOT_1445(g6751,II14825);
  not NOT_1446(g6776,g1230);
  not NOT_1447(g6777,g1346);
  not NOT_1448(g6781,g970);
  not NOT_1449(II14831,g1517);
  not NOT_1450(g6782,II14831);
  not NOT_1451(II14834,g1517);
  not NOT_1452(g6783,II14834);
  not NOT_1453(g6832,g2033);
  not NOT_1454(g6836,g1666);
  not NOT_1455(II14839,g2214);
  not NOT_1456(g6837,II14839);
  not NOT_1457(II14842,g2214);
  not NOT_1458(g6838,II14842);
  not NOT_1459(g6887,g2584);
  not NOT_1460(g6890,g2714);
  not NOT_1461(g6894,g2362);
  not NOT_1462(II14848,g2824);
  not NOT_1463(g6895,II14848);
  not NOT_1464(g6896,g2824);
  not NOT_1465(g6897,g1486);
  not NOT_1466(g6898,g2993);
  not NOT_1467(g6901,g3006);
  not NOT_1468(g6905,g3104);
  not NOT_1469(g6908,g484);
  not NOT_1470(II14857,g626);
  not NOT_1471(g6911,II14857);
  not NOT_1472(II14860,g626);
  not NOT_1473(g6912,II14860);
  not NOT_1474(g6942,g279);
  not NOT_1475(g6943,g801);
  not NOT_1476(II14865,g1237);
  not NOT_1477(g6944,II14865);
  not NOT_1478(II14868,g1237);
  not NOT_1479(g6945,II14868);
  not NOT_1480(g6974,g1151);
  not NOT_1481(g6977,g1145);
  not NOT_1482(g6978,g1245);
  not NOT_1483(II14874,g1309);
  not NOT_1484(g6979,II14874);
  not NOT_1485(II14877,g1309);
  not NOT_1486(g6980,II14877);
  not NOT_1487(g7009,g1352);
  not NOT_1488(g7013,g968);
  not NOT_1489(II14882,g1786);
  not NOT_1490(g7014,II14882);
  not NOT_1491(II14885,g1786);
  not NOT_1492(g7015,II14885);
  not NOT_1493(II14888,g1925);
  not NOT_1494(g7052,II14888);
  not NOT_1495(II14891,g1925);
  not NOT_1496(g7053,II14891);
  not NOT_1497(g7078,g1924);
  not NOT_1498(g7079,g2040);
  not NOT_1499(g7083,g1664);
  not NOT_1500(II14897,g2211);
  not NOT_1501(g7084,II14897);
  not NOT_1502(II14900,g2211);
  not NOT_1503(g7085,II14900);
  not NOT_1504(g7134,g2727);
  not NOT_1505(g7138,g2360);
  not NOT_1506(g7139,g1481);
  not NOT_1507(g7140,g2170);
  not NOT_1508(g7141,g2195);
  not NOT_1509(g7142,g8);
  not NOT_1510(g7143,g2998);
  not NOT_1511(g7146,g3013);
  not NOT_1512(g7149,g3105);
  not NOT_1513(g7152,g3136);
  not NOT_1514(g7153,g480);
  not NOT_1515(g7156,g461);
  not NOT_1516(g7157,g453);
  not NOT_1517(g7158,g1171);
  not NOT_1518(II14917,g1312);
  not NOT_1519(g7161,II14917);
  not NOT_1520(II14920,g1312);
  not NOT_1521(g7162,II14920);
  not NOT_1522(g7192,g966);
  not NOT_1523(g7193,g1491);
  not NOT_1524(II14925,g1931);
  not NOT_1525(g7194,II14925);
  not NOT_1526(II14928,g1931);
  not NOT_1527(g7195,II14928);
  not NOT_1528(g7224,g1845);
  not NOT_1529(g7227,g1839);
  not NOT_1530(g7228,g1939);
  not NOT_1531(II14934,g2003);
  not NOT_1532(g7229,II14934);
  not NOT_1533(II14937,g2003);
  not NOT_1534(g7230,II14937);
  not NOT_1535(g7259,g2046);
  not NOT_1536(g7263,g1662);
  not NOT_1537(II14942,g2480);
  not NOT_1538(g7264,II14942);
  not NOT_1539(II14945,g2480);
  not NOT_1540(g7265,II14945);
  not NOT_1541(II14948,g2619);
  not NOT_1542(g7302,II14948);
  not NOT_1543(II14951,g2619);
  not NOT_1544(g7303,II14951);
  not NOT_1545(g7328,g2618);
  not NOT_1546(g7329,g2734);
  not NOT_1547(g7333,g2358);
  not NOT_1548(II14957,g2827);
  not NOT_1549(g7334,II14957);
  not NOT_1550(g7335,g2827);
  not NOT_1551(g7336,g1476);
  not NOT_1552(g7337,g2190);
  not NOT_1553(g7338,g3002);
  not NOT_1554(g7342,g3024);
  not NOT_1555(g7345,g3139);
  not NOT_1556(g7346,g97);
  not NOT_1557(g7347,g490);
  not NOT_1558(g7348,g451);
  not NOT_1559(g7349,g1167);
  not NOT_1560(g7352,g1148);
  not NOT_1561(g7353,g1140);
  not NOT_1562(g7354,g1865);
  not NOT_1563(II14973,g2006);
  not NOT_1564(g7357,II14973);
  not NOT_1565(II14976,g2006);
  not NOT_1566(g7358,II14976);
  not NOT_1567(g7388,g1660);
  not NOT_1568(g7389,g2185);
  not NOT_1569(II14981,g2625);
  not NOT_1570(g7390,II14981);
  not NOT_1571(II14984,g2625);
  not NOT_1572(g7391,II14984);
  not NOT_1573(g7420,g2539);
  not NOT_1574(g7423,g2533);
  not NOT_1575(g7424,g2633);
  not NOT_1576(II14990,g2697);
  not NOT_1577(g7425,II14990);
  not NOT_1578(II14993,g2697);
  not NOT_1579(g7426,II14993);
  not NOT_1580(g7455,g2740);
  not NOT_1581(g7459,g2356);
  not NOT_1582(g7460,g1471);
  not NOT_1583(g7461,g2175);
  not NOT_1584(g7462,g2912);
  not NOT_1585(g7465,g2);
  not NOT_1586(g7466,g3010);
  not NOT_1587(g7471,g3036);
  not NOT_1588(g7475,g493);
  not NOT_1589(g7476,g785);
  not NOT_1590(g7477,g1177);
  not NOT_1591(g7478,g1138);
  not NOT_1592(g7479,g1861);
  not NOT_1593(g7482,g1842);
  not NOT_1594(g7483,g1834);
  not NOT_1595(g7484,g2559);
  not NOT_1596(II15012,g2700);
  not NOT_1597(g7487,II15012);
  not NOT_1598(II15015,g2700);
  not NOT_1599(g7488,II15015);
  not NOT_1600(g7518,g2354);
  not NOT_1601(II15019,g2830);
  not NOT_1602(g7519,II15019);
  not NOT_1603(g7520,g2830);
  not NOT_1604(g7521,g2200);
  not NOT_1605(g7522,g2917);
  not NOT_1606(g7527,g3018);
  not NOT_1607(g7529,g465);
  not NOT_1608(g7530,g496);
  not NOT_1609(g7531,g1180);
  not NOT_1610(g7532,g1471);
  not NOT_1611(g7533,g1871);
  not NOT_1612(g7534,g1832);
  not NOT_1613(g7535,g2555);
  not NOT_1614(g7538,g2536);
  not NOT_1615(g7539,g2528);
  not NOT_1616(g7540,g1506);
  not NOT_1617(g7541,g2180);
  not NOT_1618(g7542,g2883);
  not NOT_1619(g7545,g2920);
  not NOT_1620(g7548,g2990);
  not NOT_1621(g7549,g3028);
  not NOT_1622(g7553,g3114);
  not NOT_1623(g7554,g117);
  not NOT_1624(g7555,g1152);
  not NOT_1625(g7556,g1183);
  not NOT_1626(g7557,g1874);
  not NOT_1627(g7558,g2165);
  not NOT_1628(g7559,g2565);
  not NOT_1629(g7560,g2526);
  not NOT_1630(g7561,g1501);
  not NOT_1631(g7562,g2888);
  not NOT_1632(g7566,g2896);
  not NOT_1633(g7570,g3032);
  not NOT_1634(g7573,g3120);
  not NOT_1635(g7574,g3128);
  not NOT_1636(g7576,g468);
  not NOT_1637(g7577,g805);
  not NOT_1638(g7578,g1846);
  not NOT_1639(g7579,g1877);
  not NOT_1640(g7580,g2568);
  not NOT_1641(g7581,g1496);
  not NOT_1642(g7582,g2185);
  not NOT_1643(g7583,g2892);
  not NOT_1644(g7587,g2903);
  not NOT_1645(g7590,g1155);
  not NOT_1646(g7591,g1496);
  not NOT_1647(g7592,g2540);
  not NOT_1648(g7593,g2571);
  not NOT_1649(g7594,g2165);
  not NOT_1650(g7595,g2900);
  not NOT_1651(g7600,g2908);
  not NOT_1652(g7603,g3133);
  not NOT_1653(g7604,g471);
  not NOT_1654(g7605,g1849);
  not NOT_1655(g7606,g2190);
  not NOT_1656(g7607,g2924);
  not NOT_1657(g7610,g312);
  not NOT_1658(g7613,g1158);
  not NOT_1659(g7614,g2543);
  not NOT_1660(g7615,g3123);
  not NOT_1661(g7616,g313);
  not NOT_1662(g7619,g999);
  not NOT_1663(g7622,g1852);
  not NOT_1664(g7623,g314);
  not NOT_1665(g7626,g315);
  not NOT_1666(g7629,g403);
  not NOT_1667(g7632,g1000);
  not NOT_1668(g7635,g1693);
  not NOT_1669(g7638,g2546);
  not NOT_1670(g7639,g3094);
  not NOT_1671(g7642,g3125);
  not NOT_1672(g7643,g316);
  not NOT_1673(g7646,g318);
  not NOT_1674(g7649,g404);
  not NOT_1675(g7652,g1001);
  not NOT_1676(g7655,g1002);
  not NOT_1677(g7658,g1090);
  not NOT_1678(g7661,g1694);
  not NOT_1679(g7664,g2387);
  not NOT_1680(g7667,g3095);
  not NOT_1681(g7670,g317);
  not NOT_1682(g7673,g319);
  not NOT_1683(g7676,g402);
  not NOT_1684(g7679,g1003);
  not NOT_1685(g7682,g1005);
  not NOT_1686(g7685,g1091);
  not NOT_1687(g7688,g1695);
  not NOT_1688(g7691,g1696);
  not NOT_1689(g7694,g1784);
  not NOT_1690(g7697,g2388);
  not NOT_1691(g7700,g3096);
  not NOT_1692(g7703,g320);
  not NOT_1693(g7706,g1004);
  not NOT_1694(g7709,g1006);
  not NOT_1695(g7712,g1089);
  not NOT_1696(g7715,g1697);
  not NOT_1697(g7718,g1699);
  not NOT_1698(g7721,g1785);
  not NOT_1699(g7724,g2389);
  not NOT_1700(g7727,g2390);
  not NOT_1701(g7730,g2478);
  not NOT_1702(g7733,g1007);
  not NOT_1703(g7736,g1698);
  not NOT_1704(g7739,g1700);
  not NOT_1705(g7742,g1783);
  not NOT_1706(g7745,g2391);
  not NOT_1707(g7748,g2393);
  not NOT_1708(g7751,g2479);
  not NOT_1709(g7754,g322);
  not NOT_1710(g7757,g1701);
  not NOT_1711(g7760,g2392);
  not NOT_1712(g7763,g2394);
  not NOT_1713(g7766,g2477);
  not NOT_1714(g7769,g323);
  not NOT_1715(g7772,g659);
  not NOT_1716(g7776,g1009);
  not NOT_1717(g7779,g2395);
  not NOT_1718(g7782,g321);
  not NOT_1719(g7785,g1010);
  not NOT_1720(g7788,g1345);
  not NOT_1721(g7792,g1703);
  not NOT_1722(g7796,g1008);
  not NOT_1723(g7799,g1704);
  not NOT_1724(g7802,g2039);
  not NOT_1725(g7806,g2397);
  not NOT_1726(g7809,g1702);
  not NOT_1727(g7812,g2398);
  not NOT_1728(g7815,g2733);
  not NOT_1729(g7819,g479);
  not NOT_1730(g7822,g510);
  not NOT_1731(g7823,g2396);
  not NOT_1732(g7826,g2987);
  not NOT_1733(g7827,g478);
  not NOT_1734(g7830,g1166);
  not NOT_1735(g7833,g1196);
  not NOT_1736(g7834,g2953);
  not NOT_1737(g7837,g3044);
  not NOT_1738(g7838,g477);
  not NOT_1739(g7841,g630);
  not NOT_1740(g7842,g1165);
  not NOT_1741(g7845,g1860);
  not NOT_1742(g7848,g1890);
  not NOT_1743(g7849,g2956);
  not NOT_1744(g7852,g2981);
  not NOT_1745(g7856,g3045);
  not NOT_1746(g7857,g3055);
  not NOT_1747(g7858,g1164);
  not NOT_1748(g7861,g1316);
  not NOT_1749(g7862,g1859);
  not NOT_1750(g7865,g2554);
  not NOT_1751(g7868,g2584);
  not NOT_1752(g7869,g2959);
  not NOT_1753(g7872,g2874);
  not NOT_1754(g7877,g3046);
  not NOT_1755(g7878,g3056);
  not NOT_1756(g7879,g3065);
  not NOT_1757(g7880,g3201);
  not NOT_1758(g7888,g1858);
  not NOT_1759(g7891,g2010);
  not NOT_1760(g7892,g2553);
  not NOT_1761(g7897,g3047);
  not NOT_1762(g7898,g3057);
  not NOT_1763(g7899,g3066);
  not NOT_1764(g7900,g3075);
  not NOT_1765(II15222,g3151);
  not NOT_1766(g7901,II15222);
  not NOT_1767(g7906,g488);
  not NOT_1768(II15226,g474);
  not NOT_1769(g7909,II15226);
  not NOT_1770(g7910,g474);
  not NOT_1771(II15230,g499);
  not NOT_1772(g7911,II15230);
  not NOT_1773(g7912,g2552);
  not NOT_1774(g7915,g2704);
  not NOT_1775(g7916,g2935);
  not NOT_1776(g7919,g2963);
  not NOT_1777(g7924,g3048);
  not NOT_1778(g7925,g3058);
  not NOT_1779(g7926,g3067);
  not NOT_1780(g7927,g3076);
  not NOT_1781(g7928,g3204);
  not NOT_1782(II15256,g2950);
  not NOT_1783(g7936,II15256);
  not NOT_1784(g7949,g165);
  not NOT_1785(g7950,g142);
  not NOT_1786(g7953,g487);
  not NOT_1787(II15262,g481);
  not NOT_1788(g7956,II15262);
  not NOT_1789(g7957,g481);
  not NOT_1790(g7958,g1175);
  not NOT_1791(II15267,g1161);
  not NOT_1792(g7961,II15267);
  not NOT_1793(g7962,g1161);
  not NOT_1794(II15271,g1186);
  not NOT_1795(g7963,II15271);
  not NOT_1796(g7964,g2938);
  not NOT_1797(g7967,g2966);
  not NOT_1798(g7971,g3049);
  not NOT_1799(g7972,g3059);
  not NOT_1800(g7973,g3068);
  not NOT_1801(g7974,g3077);
  not NOT_1802(g7975,g39);
  not NOT_1803(II15288,g3109);
  not NOT_1804(g7976,II15288);
  not NOT_1805(g7989,g3191);
  not NOT_1806(g7990,g143);
  not NOT_1807(g7993,g145);
  not NOT_1808(g7996,g486);
  not NOT_1809(g7999,g485);
  not NOT_1810(g8000,g853);
  not NOT_1811(g8001,g830);
  not NOT_1812(g8004,g1174);
  not NOT_1813(II15299,g1168);
  not NOT_1814(g8007,II15299);
  not NOT_1815(g8008,g1168);
  not NOT_1816(g8009,g1869);
  not NOT_1817(II15304,g1855);
  not NOT_1818(g8012,II15304);
  not NOT_1819(g8013,g1855);
  not NOT_1820(II15308,g1880);
  not NOT_1821(g8014,II15308);
  not NOT_1822(g8015,g2941);
  not NOT_1823(g8018,g2969);
  not NOT_1824(II15313,g2930);
  not NOT_1825(g8021,II15313);
  not NOT_1826(g8022,g2930);
  not NOT_1827(II15317,g2842);
  not NOT_1828(g8023,II15317);
  not NOT_1829(g8024,g2842);
  not NOT_1830(g8025,g3050);
  not NOT_1831(g8026,g3060);
  not NOT_1832(g8027,g3069);
  not NOT_1833(g8028,g3078);
  not NOT_1834(g8029,g3083);
  not NOT_1835(II15326,g3117);
  not NOT_1836(g8030,II15326);
  not NOT_1837(II15329,g3117);
  not NOT_1838(g8031,II15329);
  not NOT_1839(g8044,g3194);
  not NOT_1840(g8045,g3207);
  not NOT_1841(g8053,g141);
  not NOT_1842(g8056,g146);
  not NOT_1843(g8059,g148);
  not NOT_1844(g8062,g169);
  not NOT_1845(g8065,g831);
  not NOT_1846(g8068,g833);
  not NOT_1847(g8071,g1173);
  not NOT_1848(g8074,g1172);
  not NOT_1849(g8075,g1547);
  not NOT_1850(g8076,g1524);
  not NOT_1851(g8079,g1868);
  not NOT_1852(II15345,g1862);
  not NOT_1853(g8082,II15345);
  not NOT_1854(g8083,g1862);
  not NOT_1855(g8084,g2563);
  not NOT_1856(II15350,g2549);
  not NOT_1857(g8087,II15350);
  not NOT_1858(g8088,g2549);
  not NOT_1859(II15354,g2574);
  not NOT_1860(g8089,II15354);
  not NOT_1861(g8090,g2944);
  not NOT_1862(g8093,g2972);
  not NOT_1863(II15359,g2858);
  not NOT_1864(g8096,II15359);
  not NOT_1865(g8097,g2858);
  not NOT_1866(g8098,g3051);
  not NOT_1867(g8099,g3061);
  not NOT_1868(g8100,g3070);
  not NOT_1869(g8101,g2997);
  not NOT_1870(g8102,g27);
  not NOT_1871(g8103,g185);
  not NOT_1872(II15369,g3129);
  not NOT_1873(g8106,II15369);
  not NOT_1874(II15372,g3129);
  not NOT_1875(g8107,II15372);
  not NOT_1876(g8120,g3197);
  not NOT_1877(g8123,g144);
  not NOT_1878(g8126,g149);
  not NOT_1879(g8129,g151);
  not NOT_1880(g8132,g170);
  not NOT_1881(g8135,g172);
  not NOT_1882(g8138,g829);
  not NOT_1883(g8141,g834);
  not NOT_1884(g8144,g836);
  not NOT_1885(g8147,g857);
  not NOT_1886(g8150,g1525);
  not NOT_1887(g8153,g1527);
  not NOT_1888(g8156,g1867);
  not NOT_1889(g8159,g1866);
  not NOT_1890(g8160,g2241);
  not NOT_1891(g8161,g2218);
  not NOT_1892(g8164,g2562);
  not NOT_1893(II15392,g2556);
  not NOT_1894(g8167,II15392);
  not NOT_1895(g8168,g2556);
  not NOT_1896(g8169,g2947);
  not NOT_1897(g8172,g2975);
  not NOT_1898(II15398,g2845);
  not NOT_1899(g8175,II15398);
  not NOT_1900(g8176,g2845);
  not NOT_1901(g8177,g3043);
  not NOT_1902(g8178,g3052);
  not NOT_1903(g8179,g3062);
  not NOT_1904(g8180,g3071);
  not NOT_1905(g8181,g48);
  not NOT_1906(g8182,g3198);
  not NOT_1907(g8183,g3188);
  not NOT_1908(g8191,g147);
  not NOT_1909(g8194,g152);
  not NOT_1910(g8197,g154);
  not NOT_1911(g8200,g168);
  not NOT_1912(g8203,g173);
  not NOT_1913(g8206,g175);
  not NOT_1914(g8209,g832);
  not NOT_1915(g8212,g837);
  not NOT_1916(g8215,g839);
  not NOT_1917(g8218,g858);
  not NOT_1918(g8221,g860);
  not NOT_1919(g8224,g1523);
  not NOT_1920(g8227,g1528);
  not NOT_1921(g8230,g1530);
  not NOT_1922(g8233,g1551);
  not NOT_1923(g8236,g2219);
  not NOT_1924(g8239,g2221);
  not NOT_1925(g8242,g2561);
  not NOT_1926(g8245,g2560);
  not NOT_1927(g8246,g2978);
  not NOT_1928(II15429,g2833);
  not NOT_1929(g8249,II15429);
  not NOT_1930(g8250,g2833);
  not NOT_1931(II15433,g2861);
  not NOT_1932(g8251,II15433);
  not NOT_1933(g8252,g2861);
  not NOT_1934(g8253,g3053);
  not NOT_1935(g8254,g3063);
  not NOT_1936(g8255,g3072);
  not NOT_1937(g8256,g30);
  not NOT_1938(g8257,g3201);
  not NOT_1939(II15442,g3235);
  not NOT_1940(g8258,II15442);
  not NOT_1941(II15445,g3236);
  not NOT_1942(g8259,II15445);
  not NOT_1943(II15448,g3237);
  not NOT_1944(g8260,II15448);
  not NOT_1945(II15451,g3238);
  not NOT_1946(g8261,II15451);
  not NOT_1947(II15454,g3239);
  not NOT_1948(g8262,II15454);
  not NOT_1949(II15457,g3240);
  not NOT_1950(g8263,II15457);
  not NOT_1951(II15460,g3241);
  not NOT_1952(g8264,II15460);
  not NOT_1953(II15463,g3242);
  not NOT_1954(g8265,II15463);
  not NOT_1955(II15466,g3243);
  not NOT_1956(g8266,II15466);
  not NOT_1957(II15469,g3244);
  not NOT_1958(g8267,II15469);
  not NOT_1959(II15472,g3245);
  not NOT_1960(g8268,II15472);
  not NOT_1961(II15475,g3246);
  not NOT_1962(g8269,II15475);
  not NOT_1963(II15478,g3247);
  not NOT_1964(g8270,II15478);
  not NOT_1965(II15481,g3248);
  not NOT_1966(g8271,II15481);
  not NOT_1967(II15484,g3249);
  not NOT_1968(g8272,II15484);
  not NOT_1969(II15487,g3250);
  not NOT_1970(g8273,II15487);
  not NOT_1971(II15490,g3251);
  not NOT_1972(g8274,II15490);
  not NOT_1973(II15493,g3252);
  not NOT_1974(g8275,II15493);
  not NOT_1975(g8276,g3253);
  not NOT_1976(g8277,g3305);
  not NOT_1977(g8278,g3337);
  not NOT_1978(II15499,g7911);
  not NOT_1979(g8284,II15499);
  not NOT_1980(g8285,g3365);
  not NOT_1981(g8286,g3461);
  not NOT_1982(g8287,g3493);
  not NOT_1983(II15505,g7963);
  not NOT_1984(g8293,II15505);
  not NOT_1985(g8294,g3521);
  not NOT_1986(g8295,g3617);
  not NOT_1987(g8296,g3649);
  not NOT_1988(II15511,g8014);
  not NOT_1989(g8302,II15511);
  not NOT_1990(g8303,g3677);
  not NOT_1991(g8304,g3773);
  not NOT_1992(g8305,g3805);
  not NOT_1993(II15517,g8089);
  not NOT_1994(g8311,II15517);
  not NOT_1995(g8312,g3833);
  not NOT_1996(g8313,g3897);
  not NOT_1997(g8317,g3919);
  not NOT_1998(II15523,g3254);
  not NOT_1999(g8321,II15523);
  not NOT_2000(II15526,g6314);
  not NOT_2001(g8324,II15526);
  not NOT_2002(II15532,g3410);
  not NOT_2003(g8330,II15532);
  not NOT_2004(II15535,g6519);
  not NOT_2005(g8333,II15535);
  not NOT_2006(II15538,g6369);
  not NOT_2007(g8336,II15538);
  not NOT_2008(II15543,g3410);
  not NOT_2009(g8341,II15543);
  not NOT_2010(II15546,g6783);
  not NOT_2011(g8344,II15546);
  not NOT_2012(II15549,g6574);
  not NOT_2013(g8347,II15549);
  not NOT_2014(II15553,g3566);
  not NOT_2015(g8351,II15553);
  not NOT_2016(II15556,g6783);
  not NOT_2017(g8354,II15556);
  not NOT_2018(II15559,g7015);
  not NOT_2019(g8357,II15559);
  not NOT_2020(II15562,g5778);
  not NOT_2021(g8360,II15562);
  not NOT_2022(II15565,g6838);
  not NOT_2023(g8363,II15565);
  not NOT_2024(II15568,g3722);
  not NOT_2025(g8366,II15568);
  not NOT_2026(II15571,g7085);
  not NOT_2027(g8369,II15571);
  not NOT_2028(II15574,g6838);
  not NOT_2029(g8372,II15574);
  not NOT_2030(II15577,g7265);
  not NOT_2031(g8375,II15577);
  not NOT_2032(II15580,g5837);
  not NOT_2033(g8378,II15580);
  not NOT_2034(II15584,g3254);
  not NOT_2035(g8382,II15584);
  not NOT_2036(II15590,g3410);
  not NOT_2037(g8388,II15590);
  not NOT_2038(II15593,g6519);
  not NOT_2039(g8391,II15593);
  not NOT_2040(II15599,g3566);
  not NOT_2041(g8397,II15599);
  not NOT_2042(II15602,g6783);
  not NOT_2043(g8400,II15602);
  not NOT_2044(II15605,g6574);
  not NOT_2045(g8403,II15605);
  not NOT_2046(II15610,g3566);
  not NOT_2047(g8408,II15610);
  not NOT_2048(II15613,g7085);
  not NOT_2049(g8411,II15613);
  not NOT_2050(II15616,g6838);
  not NOT_2051(g8414,II15616);
  not NOT_2052(II15620,g3722);
  not NOT_2053(g8418,II15620);
  not NOT_2054(II15623,g7085);
  not NOT_2055(g8421,II15623);
  not NOT_2056(II15626,g7265);
  not NOT_2057(g8424,II15626);
  not NOT_2058(II15629,g5837);
  not NOT_2059(g8427,II15629);
  not NOT_2060(II15636,g3410);
  not NOT_2061(g8434,II15636);
  not NOT_2062(II15642,g3566);
  not NOT_2063(g8440,II15642);
  not NOT_2064(II15645,g6783);
  not NOT_2065(g8443,II15645);
  not NOT_2066(II15651,g3722);
  not NOT_2067(g8449,II15651);
  not NOT_2068(II15654,g7085);
  not NOT_2069(g8452,II15654);
  not NOT_2070(II15657,g6838);
  not NOT_2071(g8455,II15657);
  not NOT_2072(II15662,g3722);
  not NOT_2073(g8460,II15662);
  not NOT_2074(II15671,g3566);
  not NOT_2075(g8469,II15671);
  not NOT_2076(II15677,g3722);
  not NOT_2077(g8475,II15677);
  not NOT_2078(II15680,g7085);
  not NOT_2079(g8478,II15680);
  not NOT_2080(II15696,g3722);
  not NOT_2081(g8494,II15696);
  not NOT_2082(g8514,g6139);
  not NOT_2083(g8530,g6156);
  not NOT_2084(g8568,g6230);
  not NOT_2085(II15771,g6000);
  not NOT_2086(g8569,II15771);
  not NOT_2087(II15779,g6000);
  not NOT_2088(g8575,II15779);
  not NOT_2089(II15784,g6000);
  not NOT_2090(g8578,II15784);
  not NOT_2091(II15787,g6000);
  not NOT_2092(g8579,II15787);
  not NOT_2093(g8580,g6281);
  not NOT_2094(g8587,g6418);
  not NOT_2095(g8594,g6623);
  not NOT_2096(II15794,g3338);
  not NOT_2097(g8602,II15794);
  not NOT_2098(g8605,g6887);
  not NOT_2099(II15800,g3494);
  not NOT_2100(g8614,II15800);
  not NOT_2101(II15803,g8107);
  not NOT_2102(g8617,II15803);
  not NOT_2103(II15806,g5550);
  not NOT_2104(g8620,II15806);
  not NOT_2105(II15810,g3338);
  not NOT_2106(g8622,II15810);
  not NOT_2107(II15815,g3650);
  not NOT_2108(g8627,II15815);
  not NOT_2109(II15818,g5596);
  not NOT_2110(g8630,II15818);
  not NOT_2111(II15822,g3494);
  not NOT_2112(g8632,II15822);
  not NOT_2113(II15827,g3806);
  not NOT_2114(g8637,II15827);
  not NOT_2115(II15830,g8031);
  not NOT_2116(g8640,II15830);
  not NOT_2117(II15833,g3338);
  not NOT_2118(g8643,II15833);
  not NOT_2119(II15836,g3366);
  not NOT_2120(g8646,II15836);
  not NOT_2121(II15839,g5613);
  not NOT_2122(g8649,II15839);
  not NOT_2123(II15843,g3650);
  not NOT_2124(g8651,II15843);
  not NOT_2125(II15847,g3878);
  not NOT_2126(g8655,II15847);
  not NOT_2127(II15850,g5627);
  not NOT_2128(g8658,II15850);
  not NOT_2129(II15853,g3494);
  not NOT_2130(g8659,II15853);
  not NOT_2131(II15856,g3522);
  not NOT_2132(g8662,II15856);
  not NOT_2133(II15859,g5638);
  not NOT_2134(g8665,II15859);
  not NOT_2135(II15863,g3806);
  not NOT_2136(g8667,II15863);
  not NOT_2137(II15866,g3878);
  not NOT_2138(g8670,II15866);
  not NOT_2139(II15869,g7976);
  not NOT_2140(g8673,II15869);
  not NOT_2141(II15873,g5655);
  not NOT_2142(g8677,II15873);
  not NOT_2143(II15876,g3650);
  not NOT_2144(g8678,II15876);
  not NOT_2145(II15879,g3678);
  not NOT_2146(g8681,II15879);
  not NOT_2147(II15882,g3878);
  not NOT_2148(g8684,II15882);
  not NOT_2149(II15887,g5693);
  not NOT_2150(g8689,II15887);
  not NOT_2151(II15890,g3806);
  not NOT_2152(g8690,II15890);
  not NOT_2153(II15893,g3834);
  not NOT_2154(g8693,II15893);
  not NOT_2155(II15896,g3878);
  not NOT_2156(g8696,II15896);
  not NOT_2157(II15899,g5626);
  not NOT_2158(g8699,II15899);
  not NOT_2159(II15902,g6486);
  not NOT_2160(g8700,II15902);
  not NOT_2161(II15909,g5745);
  not NOT_2162(g8707,II15909);
  not NOT_2163(II15912,g3878);
  not NOT_2164(g8708,II15912);
  not NOT_2165(II15915,g3878);
  not NOT_2166(g8711,II15915);
  not NOT_2167(II15918,g6643);
  not NOT_2168(g8714,II15918);
  not NOT_2169(II15922,g5654);
  not NOT_2170(g8718,II15922);
  not NOT_2171(II15925,g6751);
  not NOT_2172(g8719,II15925);
  not NOT_2173(II15932,g5423);
  not NOT_2174(g8726,II15932);
  not NOT_2175(II15935,g3878);
  not NOT_2176(g8745,II15935);
  not NOT_2177(II15938,g3338);
  not NOT_2178(g8748,II15938);
  not NOT_2179(II15942,g6945);
  not NOT_2180(g8752,II15942);
  not NOT_2181(II15946,g5692);
  not NOT_2182(g8756,II15946);
  not NOT_2183(II15949,g7053);
  not NOT_2184(g8757,II15949);
  not NOT_2185(II15955,g3878);
  not NOT_2186(g8763,II15955);
  not NOT_2187(II15958,g3878);
  not NOT_2188(g8766,II15958);
  not NOT_2189(II15961,g6051);
  not NOT_2190(g8769,II15961);
  not NOT_2191(II15964,g7554);
  not NOT_2192(g8770,II15964);
  not NOT_2193(II15967,g3494);
  not NOT_2194(g8771,II15967);
  not NOT_2195(II15971,g7195);
  not NOT_2196(g8775,II15971);
  not NOT_2197(II15975,g5744);
  not NOT_2198(g8779,II15975);
  not NOT_2199(II15978,g7303);
  not NOT_2200(g8780,II15978);
  not NOT_2201(II15983,g3878);
  not NOT_2202(g8785,II15983);
  not NOT_2203(II15986,g3878);
  not NOT_2204(g8788,II15986);
  not NOT_2205(II15989,g6053);
  not NOT_2206(g8791,II15989);
  not NOT_2207(II15992,g6055);
  not NOT_2208(g8792,II15992);
  not NOT_2209(II15995,g7577);
  not NOT_2210(g8793,II15995);
  not NOT_2211(II15998,g3650);
  not NOT_2212(g8794,II15998);
  not NOT_2213(II16002,g7391);
  not NOT_2214(g8798,II16002);
  not NOT_2215(II16006,g3878);
  not NOT_2216(g8802,II16006);
  not NOT_2217(II16009,g3878);
  not NOT_2218(g8805,II16009);
  not NOT_2219(II16012,g5390);
  not NOT_2220(g8808,II16012);
  not NOT_2221(II16015,g6056);
  not NOT_2222(g8809,II16015);
  not NOT_2223(II16018,g6058);
  not NOT_2224(g8810,II16018);
  not NOT_2225(II16021,g6060);
  not NOT_2226(g8811,II16021);
  not NOT_2227(II16024,g7591);
  not NOT_2228(g8812,II16024);
  not NOT_2229(II16027,g3806);
  not NOT_2230(g8813,II16027);
  not NOT_2231(II16031,g3878);
  not NOT_2232(g8817,II16031);
  not NOT_2233(II16034,g5396);
  not NOT_2234(g8820,II16034);
  not NOT_2235(II16037,g6061);
  not NOT_2236(g8821,II16037);
  not NOT_2237(g8822,g4602);
  not NOT_2238(II16041,g6486);
  not NOT_2239(g8823,II16041);
  not NOT_2240(II16044,g5397);
  not NOT_2241(g8824,II16044);
  not NOT_2242(II16047,g6063);
  not NOT_2243(g8825,II16047);
  not NOT_2244(II16050,g6065);
  not NOT_2245(g8826,II16050);
  not NOT_2246(II16053,g6067);
  not NOT_2247(g8827,II16053);
  not NOT_2248(II16056,g7606);
  not NOT_2249(g8828,II16056);
  not NOT_2250(II16059,g3878);
  not NOT_2251(g8829,II16059);
  not NOT_2252(II16062,g3900);
  not NOT_2253(g8832,II16062);
  not NOT_2254(II16065,g7936);
  not NOT_2255(g8835,II16065);
  not NOT_2256(II16068,g5438);
  not NOT_2257(g8836,II16068);
  not NOT_2258(II16071,g5395);
  not NOT_2259(g8839,II16071);
  not NOT_2260(II16074,g5399);
  not NOT_2261(g8840,II16074);
  not NOT_2262(II16079,g6086);
  not NOT_2263(g8843,II16079);
  not NOT_2264(II16082,g5401);
  not NOT_2265(g8844,II16082);
  not NOT_2266(II16085,g6080);
  not NOT_2267(g8845,II16085);
  not NOT_2268(g8846,g4779);
  not NOT_2269(II16089,g6751);
  not NOT_2270(g8847,II16089);
  not NOT_2271(II16092,g5402);
  not NOT_2272(g8850,II16092);
  not NOT_2273(II16095,g6082);
  not NOT_2274(g8851,II16095);
  not NOT_2275(II16098,g6084);
  not NOT_2276(g8852,II16098);
  not NOT_2277(II16101,g3878);
  not NOT_2278(g8853,II16101);
  not NOT_2279(II16104,g6448);
  not NOT_2280(g8856,II16104);
  not NOT_2281(II16107,g5398);
  not NOT_2282(g8859,II16107);
  not NOT_2283(II16110,g5404);
  not NOT_2284(g8860,II16110);
  not NOT_2285(II16114,g7936);
  not NOT_2286(g8862,II16114);
  not NOT_2287(II16117,g5473);
  not NOT_2288(g8863,II16117);
  not NOT_2289(II16120,g5400);
  not NOT_2290(g8866,II16120);
  not NOT_2291(II16123,g5406);
  not NOT_2292(g8867,II16123);
  not NOT_2293(II16128,g6103);
  not NOT_2294(g8870,II16128);
  not NOT_2295(II16131,g5408);
  not NOT_2296(g8871,II16131);
  not NOT_2297(II16134,g6099);
  not NOT_2298(g8872,II16134);
  not NOT_2299(g8873,g4955);
  not NOT_2300(II16138,g7053);
  not NOT_2301(g8874,II16138);
  not NOT_2302(II16141,g5409);
  not NOT_2303(g8877,II16141);
  not NOT_2304(II16144,g6101);
  not NOT_2305(g8878,II16144);
  not NOT_2306(II16147,g3878);
  not NOT_2307(g8879,II16147);
  not NOT_2308(II16150,g3900);
  not NOT_2309(g8882,II16150);
  not NOT_2310(II16153,g3306);
  not NOT_2311(g8885,II16153);
  not NOT_2312(II16156,g5438);
  not NOT_2313(g8888,II16156);
  not NOT_2314(II16159,g5403);
  not NOT_2315(g8891,II16159);
  not NOT_2316(II16163,g6031);
  not NOT_2317(g8893,II16163);
  not NOT_2318(II16166,g6713);
  not NOT_2319(g8894,II16166);
  not NOT_2320(II16169,g5405);
  not NOT_2321(g8897,II16169);
  not NOT_2322(II16172,g5413);
  not NOT_2323(g8898,II16172);
  not NOT_2324(II16176,g7936);
  not NOT_2325(g8900,II16176);
  not NOT_2326(II16179,g5512);
  not NOT_2327(g8901,II16179);
  not NOT_2328(II16182,g5407);
  not NOT_2329(g8904,II16182);
  not NOT_2330(II16185,g5415);
  not NOT_2331(g8905,II16185);
  not NOT_2332(II16190,g6118);
  not NOT_2333(g8908,II16190);
  not NOT_2334(II16193,g5417);
  not NOT_2335(g8909,II16193);
  not NOT_2336(II16196,g6116);
  not NOT_2337(g8910,II16196);
  not NOT_2338(g8911,g5114);
  not NOT_2339(II16200,g7303);
  not NOT_2340(g8912,II16200);
  not NOT_2341(II16203,g3878);
  not NOT_2342(g8915,II16203);
  not NOT_2343(II16206,g6448);
  not NOT_2344(g8918,II16206);
  not NOT_2345(II16209,g5438);
  not NOT_2346(g8921,II16209);
  not NOT_2347(II16212,g5411);
  not NOT_2348(g8924,II16212);
  not NOT_2349(II16215,g3462);
  not NOT_2350(g8925,II16215);
  not NOT_2351(II16218,g5473);
  not NOT_2352(g8928,II16218);
  not NOT_2353(II16221,g5412);
  not NOT_2354(g8931,II16221);
  not NOT_2355(II16225,g6042);
  not NOT_2356(g8933,II16225);
  not NOT_2357(II16228,g7015);
  not NOT_2358(g8934,II16228);
  not NOT_2359(II16231,g5414);
  not NOT_2360(g8937,II16231);
  not NOT_2361(II16234,g5420);
  not NOT_2362(g8938,II16234);
  not NOT_2363(II16238,g7936);
  not NOT_2364(g8940,II16238);
  not NOT_2365(II16241,g5556);
  not NOT_2366(g8941,II16241);
  not NOT_2367(II16244,g5416);
  not NOT_2368(g8944,II16244);
  not NOT_2369(II16247,g5422);
  not NOT_2370(g8945,II16247);
  not NOT_2371(II16252,g6134);
  not NOT_2372(g8948,II16252);
  not NOT_2373(II16255,g3900);
  not NOT_2374(g8949,II16255);
  not NOT_2375(II16258,g3306);
  not NOT_2376(g8952,II16258);
  not NOT_2377(II16261,g6448);
  not NOT_2378(g8955,II16261);
  not NOT_2379(II16264,g6713);
  not NOT_2380(g8958,II16264);
  not NOT_2381(II16267,g5473);
  not NOT_2382(g8961,II16267);
  not NOT_2383(II16270,g5418);
  not NOT_2384(g8964,II16270);
  not NOT_2385(II16273,g3618);
  not NOT_2386(g8965,II16273);
  not NOT_2387(II16276,g5512);
  not NOT_2388(g8968,II16276);
  not NOT_2389(II16279,g5419);
  not NOT_2390(g8971,II16279);
  not NOT_2391(II16283,g6046);
  not NOT_2392(g8973,II16283);
  not NOT_2393(II16286,g7265);
  not NOT_2394(g8974,II16286);
  not NOT_2395(II16289,g5421);
  not NOT_2396(g8977,II16289);
  not NOT_2397(II16292,g5426);
  not NOT_2398(g8978,II16292);
  not NOT_2399(II16296,g3306);
  not NOT_2400(g8980,II16296);
  not NOT_2401(g8983,g6486);
  not NOT_2402(II16300,g3462);
  not NOT_2403(g8984,II16300);
  not NOT_2404(II16303,g6713);
  not NOT_2405(g8987,II16303);
  not NOT_2406(II16306,g7015);
  not NOT_2407(g8990,II16306);
  not NOT_2408(II16309,g5512);
  not NOT_2409(g8993,II16309);
  not NOT_2410(II16312,g5424);
  not NOT_2411(g8996,II16312);
  not NOT_2412(II16315,g3774);
  not NOT_2413(g8997,II16315);
  not NOT_2414(II16318,g5556);
  not NOT_2415(g9000,II16318);
  not NOT_2416(II16321,g5425);
  not NOT_2417(g9003,II16321);
  not NOT_2418(II16325,g6052);
  not NOT_2419(g9005,II16325);
  not NOT_2420(II16328,g3900);
  not NOT_2421(g9006,II16328);
  not NOT_2422(II16332,g3462);
  not NOT_2423(g9010,II16332);
  not NOT_2424(II16335,g3618);
  not NOT_2425(g9013,II16335);
  not NOT_2426(II16338,g7015);
  not NOT_2427(g9016,II16338);
  not NOT_2428(II16341,g7265);
  not NOT_2429(g9019,II16341);
  not NOT_2430(II16344,g5556);
  not NOT_2431(g9022,II16344);
  not NOT_2432(II16347,g5427);
  not NOT_2433(g9025,II16347);
  not NOT_2434(g9027,g5679);
  not NOT_2435(II16354,g3618);
  not NOT_2436(g9035,II16354);
  not NOT_2437(II16357,g3774);
  not NOT_2438(g9038,II16357);
  not NOT_2439(II16360,g7265);
  not NOT_2440(g9041,II16360);
  not NOT_2441(II16363,g3900);
  not NOT_2442(g9044,II16363);
  not NOT_2443(g9050,g5731);
  not NOT_2444(II16372,g3774);
  not NOT_2445(g9058,II16372);
  not NOT_2446(g9067,g5789);
  not NOT_2447(g9084,g5848);
  not NOT_2448(II16432,g3366);
  not NOT_2449(g9128,II16432);
  not NOT_2450(II16438,g3522);
  not NOT_2451(g9134,II16438);
  not NOT_2452(II16444,g3678);
  not NOT_2453(g9140,II16444);
  not NOT_2454(II16450,g3834);
  not NOT_2455(g9146,II16450);
  not NOT_2456(II16453,g7936);
  not NOT_2457(g9149,II16453);
  not NOT_2458(g9150,g5893);
  not NOT_2459(II16457,g7936);
  not NOT_2460(g9159,II16457);
  not NOT_2461(g9160,g6170);
  not NOT_2462(g9161,g5852);
  not NOT_2463(II16462,g5438);
  not NOT_2464(g9170,II16462);
  not NOT_2465(II16465,g6000);
  not NOT_2466(g9173,II16465);
  not NOT_2467(g9174,g5932);
  not NOT_2468(II16469,g7936);
  not NOT_2469(g9183,II16469);
  not NOT_2470(II16472,g7901);
  not NOT_2471(g9184,II16472);
  not NOT_2472(g9187,g5803);
  not NOT_2473(II16476,g6448);
  not NOT_2474(g9196,II16476);
  not NOT_2475(II16479,g5438);
  not NOT_2476(g9199,II16479);
  not NOT_2477(II16482,g6000);
  not NOT_2478(g9202,II16482);
  not NOT_2479(g9203,g5899);
  not NOT_2480(II16486,g5473);
  not NOT_2481(g9212,II16486);
  not NOT_2482(II16489,g6000);
  not NOT_2483(g9215,II16489);
  not NOT_2484(g9216,g5966);
  not NOT_2485(II16493,g7936);
  not NOT_2486(g9225,II16493);
  not NOT_2487(g9226,g5434);
  not NOT_2488(g9227,g5587);
  not NOT_2489(g9228,g7667);
  not NOT_2490(II16499,g7901);
  not NOT_2491(g9229,II16499);
  not NOT_2492(g9232,g5752);
  not NOT_2493(II16504,g3306);
  not NOT_2494(g9242,II16504);
  not NOT_2495(II16507,g6448);
  not NOT_2496(g9245,II16507);
  not NOT_2497(g9248,g5859);
  not NOT_2498(II16511,g6713);
  not NOT_2499(g9257,II16511);
  not NOT_2500(II16514,g5473);
  not NOT_2501(g9260,II16514);
  not NOT_2502(II16517,g6000);
  not NOT_2503(g9263,II16517);
  not NOT_2504(g9264,g5938);
  not NOT_2505(II16521,g5512);
  not NOT_2506(g9273,II16521);
  not NOT_2507(II16524,g6000);
  not NOT_2508(g9276,II16524);
  not NOT_2509(g9277,g5995);
  not NOT_2510(g9286,g6197);
  not NOT_2511(g9287,g6638);
  not NOT_2512(g9288,g5363);
  not NOT_2513(g9289,g5379);
  not NOT_2514(II16532,g7901);
  not NOT_2515(g9290,II16532);
  not NOT_2516(g9293,g5703);
  not NOT_2517(II16538,g3306);
  not NOT_2518(g9303,II16538);
  not NOT_2519(II16541,g5438);
  not NOT_2520(g9306,II16541);
  not NOT_2521(II16544,g6054);
  not NOT_2522(g9309,II16544);
  not NOT_2523(g9310,g5811);
  not NOT_2524(II16549,g3462);
  not NOT_2525(g9320,II16549);
  not NOT_2526(II16552,g6713);
  not NOT_2527(g9323,II16552);
  not NOT_2528(g9326,g5906);
  not NOT_2529(II16556,g7015);
  not NOT_2530(g9335,II16556);
  not NOT_2531(II16559,g5512);
  not NOT_2532(g9338,II16559);
  not NOT_2533(II16562,g6000);
  not NOT_2534(g9341,II16562);
  not NOT_2535(g9342,g5972);
  not NOT_2536(II16566,g5556);
  not NOT_2537(g9351,II16566);
  not NOT_2538(II16569,g6000);
  not NOT_2539(g9354,II16569);
  not NOT_2540(g9355,g7639);
  not NOT_2541(g9356,g5665);
  not NOT_2542(II16578,g6448);
  not NOT_2543(g9368,II16578);
  not NOT_2544(II16581,g5438);
  not NOT_2545(g9371,II16581);
  not NOT_2546(g9374,g5761);
  not NOT_2547(II16587,g3462);
  not NOT_2548(g9384,II16587);
  not NOT_2549(II16590,g5473);
  not NOT_2550(g9387,II16590);
  not NOT_2551(II16593,g6059);
  not NOT_2552(g9390,II16593);
  not NOT_2553(g9391,g5867);
  not NOT_2554(II16598,g3618);
  not NOT_2555(g9401,II16598);
  not NOT_2556(II16601,g7015);
  not NOT_2557(g9404,II16601);
  not NOT_2558(g9407,g5945);
  not NOT_2559(II16605,g7265);
  not NOT_2560(g9416,II16605);
  not NOT_2561(II16608,g5556);
  not NOT_2562(g9419,II16608);
  not NOT_2563(II16611,g6000);
  not NOT_2564(g9422,II16611);
  not NOT_2565(g9423,g5428);
  not NOT_2566(g9424,g5469);
  not NOT_2567(g9425,g5346);
  not NOT_2568(g9426,g5543);
  not NOT_2569(g9427,g5645);
  not NOT_2570(II16624,g3306);
  not NOT_2571(g9443,II16624);
  not NOT_2572(II16627,g6448);
  not NOT_2573(g9446,II16627);
  not NOT_2574(II16630,g6057);
  not NOT_2575(g9449,II16630);
  not NOT_2576(II16633,g6486);
  not NOT_2577(g9450,II16633);
  not NOT_2578(g9453,g5717);
  not NOT_2579(II16641,g6713);
  not NOT_2580(g9465,II16641);
  not NOT_2581(II16644,g5473);
  not NOT_2582(g9468,II16644);
  not NOT_2583(g9471,g5820);
  not NOT_2584(II16650,g3618);
  not NOT_2585(g9481,II16650);
  not NOT_2586(II16653,g5512);
  not NOT_2587(g9484,II16653);
  not NOT_2588(II16656,g6066);
  not NOT_2589(g9487,II16656);
  not NOT_2590(g9488,g5914);
  not NOT_2591(II16661,g3774);
  not NOT_2592(g9498,II16661);
  not NOT_2593(II16664,g7265);
  not NOT_2594(g9501,II16664);
  not NOT_2595(g9504,g6149);
  not NOT_2596(g9505,g6227);
  not NOT_2597(g9506,g6444);
  not NOT_2598(g9507,g5953);
  not NOT_2599(II16677,g3306);
  not NOT_2600(g9524,II16677);
  not NOT_2601(g9527,g5508);
  not NOT_2602(II16681,g6643);
  not NOT_2603(g9528,II16681);
  not NOT_2604(II16684,g6486);
  not NOT_2605(g9531,II16684);
  not NOT_2606(g9569,g5683);
  not NOT_2607(II16694,g3462);
  not NOT_2608(g9585,II16694);
  not NOT_2609(II16697,g6713);
  not NOT_2610(g9588,II16697);
  not NOT_2611(II16700,g6064);
  not NOT_2612(g9591,II16700);
  not NOT_2613(II16703,g6751);
  not NOT_2614(g9592,II16703);
  not NOT_2615(g9595,g5775);
  not NOT_2616(II16711,g7015);
  not NOT_2617(g9607,II16711);
  not NOT_2618(II16714,g5512);
  not NOT_2619(g9610,II16714);
  not NOT_2620(g9613,g5876);
  not NOT_2621(II16720,g3774);
  not NOT_2622(g9623,II16720);
  not NOT_2623(II16723,g5556);
  not NOT_2624(g9626,II16723);
  not NOT_2625(II16726,g6085);
  not NOT_2626(g9629,II16726);
  not NOT_2627(II16741,g6062);
  not NOT_2628(g9640,II16741);
  not NOT_2629(II16744,g3338);
  not NOT_2630(g9641,II16744);
  not NOT_2631(II16747,g6643);
  not NOT_2632(g9644,II16747);
  not NOT_2633(g9649,g5982);
  not NOT_2634(II16759,g3462);
  not NOT_2635(g9666,II16759);
  not NOT_2636(g9669,g5552);
  not NOT_2637(II16763,g6945);
  not NOT_2638(g9670,II16763);
  not NOT_2639(II16766,g6751);
  not NOT_2640(g9673,II16766);
  not NOT_2641(g9711,g5735);
  not NOT_2642(II16776,g3618);
  not NOT_2643(g9727,II16776);
  not NOT_2644(II16779,g7015);
  not NOT_2645(g9730,II16779);
  not NOT_2646(II16782,g6083);
  not NOT_2647(g9733,II16782);
  not NOT_2648(II16785,g7053);
  not NOT_2649(g9734,II16785);
  not NOT_2650(g9737,g5834);
  not NOT_2651(II16793,g7265);
  not NOT_2652(g9749,II16793);
  not NOT_2653(II16796,g5556);
  not NOT_2654(g9752,II16796);
  not NOT_2655(g9755,g5431);
  not NOT_2656(g9756,g5504);
  not NOT_2657(g9757,g5601);
  not NOT_2658(g9758,g5618);
  not NOT_2659(II16811,g3338);
  not NOT_2660(g9767,II16811);
  not NOT_2661(II16814,g6486);
  not NOT_2662(g9770,II16814);
  not NOT_2663(II16832,g6081);
  not NOT_2664(g9786,II16832);
  not NOT_2665(II16835,g3494);
  not NOT_2666(g9787,II16835);
  not NOT_2667(II16838,g6945);
  not NOT_2668(g9790,II16838);
  not NOT_2669(g9795,g6019);
  not NOT_2670(II16850,g3618);
  not NOT_2671(g9812,II16850);
  not NOT_2672(g9815,g5598);
  not NOT_2673(II16854,g7195);
  not NOT_2674(g9816,II16854);
  not NOT_2675(II16857,g7053);
  not NOT_2676(g9819,II16857);
  not NOT_2677(g9857,g5793);
  not NOT_2678(II16867,g3774);
  not NOT_2679(g9873,II16867);
  not NOT_2680(II16870,g7265);
  not NOT_2681(g9876,II16870);
  not NOT_2682(II16873,g6102);
  not NOT_2683(g9879,II16873);
  not NOT_2684(II16876,g7303);
  not NOT_2685(g9880,II16876);
  not NOT_2686(g9884,g6310);
  not NOT_2687(g9885,g6905);
  not NOT_2688(g9886,g7149);
  not NOT_2689(II16897,g6643);
  not NOT_2690(g9895,II16897);
  not NOT_2691(II16900,g6486);
  not NOT_2692(g9898,II16900);
  not NOT_2693(II16915,g3494);
  not NOT_2694(g9913,II16915);
  not NOT_2695(II16918,g6751);
  not NOT_2696(g9916,II16918);
  not NOT_2697(II16936,g6100);
  not NOT_2698(g9932,II16936);
  not NOT_2699(II16939,g3650);
  not NOT_2700(g9933,II16939);
  not NOT_2701(II16942,g7195);
  not NOT_2702(g9936,II16942);
  not NOT_2703(g9941,g6035);
  not NOT_2704(II16954,g3774);
  not NOT_2705(g9958,II16954);
  not NOT_2706(g9961,g5615);
  not NOT_2707(II16958,g7391);
  not NOT_2708(g9962,II16958);
  not NOT_2709(II16961,g7303);
  not NOT_2710(g9965,II16961);
  not NOT_2711(II16972,g3900);
  not NOT_2712(g10004,II16972);
  not NOT_2713(g10015,g5292);
  not NOT_2714(II16984,g7936);
  not NOT_2715(g10016,II16984);
  not NOT_2716(II16987,g6079);
  not NOT_2717(g10017,II16987);
  not NOT_2718(II16990,g3338);
  not NOT_2719(g10018,II16990);
  not NOT_2720(II16993,g6643);
  not NOT_2721(g10021,II16993);
  not NOT_2722(II17009,g6945);
  not NOT_2723(g10049,II17009);
  not NOT_2724(II17012,g6751);
  not NOT_2725(g10052,II17012);
  not NOT_2726(II17027,g3650);
  not NOT_2727(g10067,II17027);
  not NOT_2728(II17030,g7053);
  not NOT_2729(g10070,II17030);
  not NOT_2730(II17048,g6117);
  not NOT_2731(g10086,II17048);
  not NOT_2732(II17051,g3806);
  not NOT_2733(g10087,II17051);
  not NOT_2734(II17054,g7391);
  not NOT_2735(g10090,II17054);
  not NOT_2736(II17066,g3900);
  not NOT_2737(g10096,II17066);
  not NOT_2738(g10099,g7700);
  not NOT_2739(II17070,g7528);
  not NOT_2740(g10100,II17070);
  not NOT_2741(II17081,g3338);
  not NOT_2742(g10109,II17081);
  not NOT_2743(g10124,g5326);
  not NOT_2744(II17097,g7936);
  not NOT_2745(g10125,II17097);
  not NOT_2746(II17100,g6098);
  not NOT_2747(g10126,II17100);
  not NOT_2748(II17103,g3494);
  not NOT_2749(g10127,II17103);
  not NOT_2750(II17106,g6945);
  not NOT_2751(g10130,II17106);
  not NOT_2752(II17122,g7195);
  not NOT_2753(g10158,II17122);
  not NOT_2754(II17125,g7053);
  not NOT_2755(g10161,II17125);
  not NOT_2756(II17140,g3806);
  not NOT_2757(g10176,II17140);
  not NOT_2758(II17143,g7303);
  not NOT_2759(g10179,II17143);
  not NOT_2760(II17159,g3900);
  not NOT_2761(g10189,II17159);
  not NOT_2762(II17184,g3494);
  not NOT_2763(g10214,II17184);
  not NOT_2764(g10229,g5349);
  not NOT_2765(II17200,g7936);
  not NOT_2766(g10230,II17200);
  not NOT_2767(II17203,g6115);
  not NOT_2768(g10231,II17203);
  not NOT_2769(II17206,g3650);
  not NOT_2770(g10232,II17206);
  not NOT_2771(II17209,g7195);
  not NOT_2772(g10235,II17209);
  not NOT_2773(II17225,g7391);
  not NOT_2774(g10263,II17225);
  not NOT_2775(II17228,g7303);
  not NOT_2776(g10266,II17228);
  not NOT_2777(II17235,g3900);
  not NOT_2778(g10273,II17235);
  not NOT_2779(II17238,g3900);
  not NOT_2780(g10276,II17238);
  not NOT_2781(II17278,g3650);
  not NOT_2782(g10316,II17278);
  not NOT_2783(g10331,g5366);
  not NOT_2784(II17294,g7936);
  not NOT_2785(g10332,II17294);
  not NOT_2786(II17297,g6130);
  not NOT_2787(g10333,II17297);
  not NOT_2788(II17300,g3806);
  not NOT_2789(g10334,II17300);
  not NOT_2790(II17303,g7391);
  not NOT_2791(g10337,II17303);
  not NOT_2792(II17311,g3900);
  not NOT_2793(g10357,II17311);
  not NOT_2794(II17363,g3806);
  not NOT_2795(g10409,II17363);
  not NOT_2796(II17370,g3900);
  not NOT_2797(g10416,II17370);
  not NOT_2798(II17373,g3900);
  not NOT_2799(g10419,II17373);
  not NOT_2800(g10424,g7910);
  not NOT_2801(g10481,g7826);
  not NOT_2802(II17433,g3900);
  not NOT_2803(g10482,II17433);
  not NOT_2804(g10486,g7957);
  not NOT_2805(g10500,g7962);
  not NOT_2806(II17483,g3900);
  not NOT_2807(g10542,II17483);
  not NOT_2808(II17486,g3900);
  not NOT_2809(g10545,II17486);
  not NOT_2810(g10549,g7999);
  not NOT_2811(g10560,g8008);
  not NOT_2812(g10574,g8013);
  not NOT_2813(II17527,g3900);
  not NOT_2814(g10601,II17527);
  not NOT_2815(g10606,g8074);
  not NOT_2816(g10617,g8083);
  not NOT_2817(g10631,g8088);
  not NOT_2818(II17557,g3900);
  not NOT_2819(g10646,II17557);
  not NOT_2820(g10653,g8159);
  not NOT_2821(g10664,g8168);
  not NOT_2822(g10683,g8245);
  not NOT_2823(g10694,g4326);
  not NOT_2824(g10714,g4495);
  not NOT_2825(g10730,g6173);
  not NOT_2826(g10735,g4671);
  not NOT_2827(g10749,g6205);
  not NOT_2828(g10754,g4848);
  not NOT_2829(g10765,g6048);
  not NOT_2830(g10766,g6676);
  not NOT_2831(g10767,g6294);
  not NOT_2832(g10772,g6978);
  not NOT_2833(g10773,g6431);
  not NOT_2834(II17627,g7575);
  not NOT_2835(g10779,II17627);
  not NOT_2836(g10783,g7228);
  not NOT_2837(II17632,g6183);
  not NOT_2838(g10787,II17632);
  not NOT_2839(g10788,g7424);
  not NOT_2840(II17637,g6204);
  not NOT_2841(g10792,II17637);
  not NOT_2842(II17641,g6215);
  not NOT_2843(g10796,II17641);
  not NOT_2844(II17645,g6288);
  not NOT_2845(g10800,II17645);
  not NOT_2846(II17649,g6293);
  not NOT_2847(g10804,II17649);
  not NOT_2848(II17653,g6304);
  not NOT_2849(g10808,II17653);
  not NOT_2850(g10809,g5701);
  not NOT_2851(II17658,g6367);
  not NOT_2852(g10813,II17658);
  not NOT_2853(II17662,g6425);
  not NOT_2854(g10817,II17662);
  not NOT_2855(II17666,g6430);
  not NOT_2856(g10821,II17666);
  not NOT_2857(II17670,g6441);
  not NOT_2858(g10825,II17670);
  not NOT_2859(II17673,g8107);
  not NOT_2860(g10826,II17673);
  not NOT_2861(g10829,g5749);
  not NOT_2862(II17677,g6517);
  not NOT_2863(g10830,II17677);
  not NOT_2864(II17681,g6572);
  not NOT_2865(g10834,II17681);
  not NOT_2866(II17685,g6630);
  not NOT_2867(g10838,II17685);
  not NOT_2868(II17689,g6635);
  not NOT_2869(g10842,II17689);
  not NOT_2870(II17692,g8107);
  not NOT_2871(g10843,II17692);
  not NOT_2872(g10846,g5799);
  not NOT_2873(g10847,g5800);
  not NOT_2874(g10848,g5801);
  not NOT_2875(II17698,g6711);
  not NOT_2876(g10849,II17698);
  not NOT_2877(II17701,g6781);
  not NOT_2878(g10850,II17701);
  not NOT_2879(II17705,g6836);
  not NOT_2880(g10854,II17705);
  not NOT_2881(II17709,g6894);
  not NOT_2882(g10858,II17709);
  not NOT_2883(II17712,g8031);
  not NOT_2884(g10859,II17712);
  not NOT_2885(II17715,g8107);
  not NOT_2886(g10862,II17715);
  not NOT_2887(g10865,g6131);
  not NOT_2888(g10866,g5849);
  not NOT_2889(g10867,g5850);
  not NOT_2890(II17721,g6641);
  not NOT_2891(g10868,II17721);
  not NOT_2892(II17724,g6942);
  not NOT_2893(g10869,II17724);
  not NOT_2894(II17727,g7013);
  not NOT_2895(g10870,II17727);
  not NOT_2896(II17730,g7083);
  not NOT_2897(g10871,II17730);
  not NOT_2898(II17734,g7138);
  not NOT_2899(g10875,II17734);
  not NOT_2900(II17737,g6000);
  not NOT_2901(g10876,II17737);
  not NOT_2902(II17740,g8031);
  not NOT_2903(g10877,II17740);
  not NOT_2904(II17743,g8107);
  not NOT_2905(g10880,II17743);
  not NOT_2906(II17746,g8107);
  not NOT_2907(g10883,II17746);
  not NOT_2908(g10886,g5889);
  not NOT_2909(II17750,g7157);
  not NOT_2910(g10887,II17750);
  not NOT_2911(II17753,g6943);
  not NOT_2912(g10888,II17753);
  not NOT_2913(II17756,g7192);
  not NOT_2914(g10889,II17756);
  not NOT_2915(II17759,g7263);
  not NOT_2916(g10890,II17759);
  not NOT_2917(II17762,g7333);
  not NOT_2918(g10891,II17762);
  not NOT_2919(II17765,g7976);
  not NOT_2920(g10892,II17765);
  not NOT_2921(II17768,g8031);
  not NOT_2922(g10895,II17768);
  not NOT_2923(II17771,g8107);
  not NOT_2924(g10898,II17771);
  not NOT_2925(II17774,g8107);
  not NOT_2926(g10901,II17774);
  not NOT_2927(g10904,g5922);
  not NOT_2928(g10905,g5923);
  not NOT_2929(g10906,g5924);
  not NOT_2930(II17780,g7348);
  not NOT_2931(g10907,II17780);
  not NOT_2932(II17783,g7353);
  not NOT_2933(g10908,II17783);
  not NOT_2934(II17786,g7193);
  not NOT_2935(g10909,II17786);
  not NOT_2936(II17789,g7388);
  not NOT_2937(g10910,II17789);
  not NOT_2938(II17792,g7459);
  not NOT_2939(g10911,II17792);
  not NOT_2940(II17795,g7976);
  not NOT_2941(g10912,II17795);
  not NOT_2942(II17798,g8031);
  not NOT_2943(g10915,II17798);
  not NOT_2944(II17801,g8107);
  not NOT_2945(g10918,II17801);
  not NOT_2946(II17804,g8031);
  not NOT_2947(g10921,II17804);
  not NOT_2948(II17807,g8107);
  not NOT_2949(g10924,II17807);
  not NOT_2950(g10927,g6153);
  not NOT_2951(g10928,g5951);
  not NOT_2952(g10929,g5952);
  not NOT_2953(II17813,g5707);
  not NOT_2954(g10930,II17813);
  not NOT_2955(II17816,g7346);
  not NOT_2956(g10931,II17816);
  not NOT_2957(II17819,g6448);
  not NOT_2958(g10932,II17819);
  not NOT_2959(II17822,g7478);
  not NOT_2960(g10933,II17822);
  not NOT_2961(II17825,g7483);
  not NOT_2962(g10934,II17825);
  not NOT_2963(II17828,g7389);
  not NOT_2964(g10935,II17828);
  not NOT_2965(II17831,g7518);
  not NOT_2966(g10936,II17831);
  not NOT_2967(II17834,g7976);
  not NOT_2968(g10937,II17834);
  not NOT_2969(II17837,g8031);
  not NOT_2970(g10940,II17837);
  not NOT_2971(II17840,g8107);
  not NOT_2972(g10943,II17840);
  not NOT_2973(II17843,g8031);
  not NOT_2974(g10946,II17843);
  not NOT_2975(II17846,g8107);
  not NOT_2976(g10949,II17846);
  not NOT_2977(II17849,g8103);
  not NOT_2978(g10952,II17849);
  not NOT_2979(g10961,g5978);
  not NOT_2980(g10962,g5979);
  not NOT_2981(II17854,g6232);
  not NOT_2982(g10963,II17854);
  not NOT_2983(II17857,g6448);
  not NOT_2984(g10966,II17857);
  not NOT_2985(II17860,g5765);
  not NOT_2986(g10967,II17860);
  not NOT_2987(II17863,g7476);
  not NOT_2988(g10968,II17863);
  not NOT_2989(II17866,g6713);
  not NOT_2990(g10969,II17866);
  not NOT_2991(II17869,g7534);
  not NOT_2992(g10972,II17869);
  not NOT_2993(II17872,g7539);
  not NOT_2994(g10973,II17872);
  not NOT_2995(II17875,g7976);
  not NOT_2996(g10974,II17875);
  not NOT_2997(II17878,g8031);
  not NOT_2998(g10977,II17878);
  not NOT_2999(II17881,g7976);
  not NOT_3000(g10980,II17881);
  not NOT_3001(II17884,g8031);
  not NOT_3002(g10983,II17884);
  not NOT_3003(g10986,g6014);
  not NOT_3004(g10987,g6015);
  not NOT_3005(II17889,g6314);
  not NOT_3006(g10988,II17889);
  not NOT_3007(II17892,g6232);
  not NOT_3008(g10991,II17892);
  not NOT_3009(II17895,g6448);
  not NOT_3010(g10994,II17895);
  not NOT_3011(II17898,g6643);
  not NOT_3012(g10995,II17898);
  not NOT_3013(II17901,g6369);
  not NOT_3014(g10996,II17901);
  not NOT_3015(II17904,g6713);
  not NOT_3016(g10999,II17904);
  not NOT_3017(II17907,g5824);
  not NOT_3018(g11002,II17907);
  not NOT_3019(II17910,g7532);
  not NOT_3020(g11003,II17910);
  not NOT_3021(II17913,g7015);
  not NOT_3022(g11004,II17913);
  not NOT_3023(II17916,g7560);
  not NOT_3024(g11007,II17916);
  not NOT_3025(II17919,g7976);
  not NOT_3026(g11008,II17919);
  not NOT_3027(II17922,g8031);
  not NOT_3028(g11011,II17922);
  not NOT_3029(II17925,g7976);
  not NOT_3030(g11014,II17925);
  not NOT_3031(II17928,g8031);
  not NOT_3032(g11017,II17928);
  not NOT_3033(g11020,g6029);
  not NOT_3034(g11021,g6030);
  not NOT_3035(II17933,g3254);
  not NOT_3036(g11022,II17933);
  not NOT_3037(II17936,g6314);
  not NOT_3038(g11025,II17936);
  not NOT_3039(II17939,g6232);
  not NOT_3040(g11028,II17939);
  not NOT_3041(II17942,g5548);
  not NOT_3042(g11031,II17942);
  not NOT_3043(II17945,g5668);
  not NOT_3044(g11032,II17945);
  not NOT_3045(II17948,g6643);
  not NOT_3046(g11035,II17948);
  not NOT_3047(II17951,g6519);
  not NOT_3048(g11036,II17951);
  not NOT_3049(II17954,g6369);
  not NOT_3050(g11039,II17954);
  not NOT_3051(II17957,g6713);
  not NOT_3052(g11042,II17957);
  not NOT_3053(II17960,g6945);
  not NOT_3054(g11045,II17960);
  not NOT_3055(II17963,g6574);
  not NOT_3056(g11048,II17963);
  not NOT_3057(II17966,g7015);
  not NOT_3058(g11051,II17966);
  not NOT_3059(II17969,g5880);
  not NOT_3060(g11054,II17969);
  not NOT_3061(II17972,g7558);
  not NOT_3062(g11055,II17972);
  not NOT_3063(II17975,g7265);
  not NOT_3064(g11056,II17975);
  not NOT_3065(II17978,g7795);
  not NOT_3066(g11059,II17978);
  not NOT_3067(II17981,g7976);
  not NOT_3068(g11063,II17981);
  not NOT_3069(II17984,g7976);
  not NOT_3070(g11066,II17984);
  not NOT_3071(g11069,g8257);
  not NOT_3072(g11078,g6041);
  not NOT_3073(II17989,g3254);
  not NOT_3074(g11079,II17989);
  not NOT_3075(II17992,g6314);
  not NOT_3076(g11082,II17992);
  not NOT_3077(II17995,g6232);
  not NOT_3078(g11085,II17995);
  not NOT_3079(II17998,g5668);
  not NOT_3080(g11088,II17998);
  not NOT_3081(II18001,g6643);
  not NOT_3082(g11091,II18001);
  not NOT_3083(II18004,g3410);
  not NOT_3084(g11092,II18004);
  not NOT_3085(II18007,g6519);
  not NOT_3086(g11095,II18007);
  not NOT_3087(II18010,g6369);
  not NOT_3088(g11098,II18010);
  not NOT_3089(II18013,g5594);
  not NOT_3090(g11101,II18013);
  not NOT_3091(II18016,g5720);
  not NOT_3092(g11102,II18016);
  not NOT_3093(II18019,g6945);
  not NOT_3094(g11105,II18019);
  not NOT_3095(II18022,g6783);
  not NOT_3096(g11108,II18022);
  not NOT_3097(II18025,g6574);
  not NOT_3098(g11111,II18025);
  not NOT_3099(II18028,g7015);
  not NOT_3100(g11114,II18028);
  not NOT_3101(II18031,g7195);
  not NOT_3102(g11117,II18031);
  not NOT_3103(II18034,g6838);
  not NOT_3104(g11120,II18034);
  not NOT_3105(II18037,g7265);
  not NOT_3106(g11123,II18037);
  not NOT_3107(II18040,g7976);
  not NOT_3108(g11126,II18040);
  not NOT_3109(II18043,g7976);
  not NOT_3110(g11129,II18043);
  not NOT_3111(II18046,g3254);
  not NOT_3112(g11132,II18046);
  not NOT_3113(II18049,g6314);
  not NOT_3114(g11135,II18049);
  not NOT_3115(II18052,g6232);
  not NOT_3116(g11138,II18052);
  not NOT_3117(II18055,g5668);
  not NOT_3118(g11141,II18055);
  not NOT_3119(II18058,g6643);
  not NOT_3120(g11144,II18058);
  not NOT_3121(II18061,g3410);
  not NOT_3122(g11145,II18061);
  not NOT_3123(II18064,g6519);
  not NOT_3124(g11148,II18064);
  not NOT_3125(II18067,g6369);
  not NOT_3126(g11151,II18067);
  not NOT_3127(II18070,g5720);
  not NOT_3128(g11154,II18070);
  not NOT_3129(II18073,g6945);
  not NOT_3130(g11157,II18073);
  not NOT_3131(II18076,g3566);
  not NOT_3132(g11160,II18076);
  not NOT_3133(II18079,g6783);
  not NOT_3134(g11163,II18079);
  not NOT_3135(II18082,g6574);
  not NOT_3136(g11166,II18082);
  not NOT_3137(II18085,g5611);
  not NOT_3138(g11169,II18085);
  not NOT_3139(II18088,g5778);
  not NOT_3140(g11170,II18088);
  not NOT_3141(II18091,g7195);
  not NOT_3142(g11173,II18091);
  not NOT_3143(II18094,g7085);
  not NOT_3144(g11176,II18094);
  not NOT_3145(II18097,g6838);
  not NOT_3146(g11179,II18097);
  not NOT_3147(II18100,g7265);
  not NOT_3148(g11182,II18100);
  not NOT_3149(II18103,g7391);
  not NOT_3150(g11185,II18103);
  not NOT_3151(g11190,g3999);
  not NOT_3152(II18121,g3254);
  not NOT_3153(g11199,II18121);
  not NOT_3154(II18124,g6314);
  not NOT_3155(g11202,II18124);
  not NOT_3156(II18127,g6232);
  not NOT_3157(g11205,II18127);
  not NOT_3158(II18130,g5547);
  not NOT_3159(g11208,II18130);
  not NOT_3160(II18133,g6448);
  not NOT_3161(g11209,II18133);
  not NOT_3162(II18136,g5668);
  not NOT_3163(g11210,II18136);
  not NOT_3164(II18139,g6643);
  not NOT_3165(g11213,II18139);
  not NOT_3166(II18142,g3410);
  not NOT_3167(g11216,II18142);
  not NOT_3168(II18145,g6519);
  not NOT_3169(g11219,II18145);
  not NOT_3170(II18148,g6369);
  not NOT_3171(g11222,II18148);
  not NOT_3172(II18151,g5720);
  not NOT_3173(g11225,II18151);
  not NOT_3174(II18154,g6945);
  not NOT_3175(g11228,II18154);
  not NOT_3176(II18157,g3566);
  not NOT_3177(g11231,II18157);
  not NOT_3178(II18160,g6783);
  not NOT_3179(g11234,II18160);
  not NOT_3180(II18163,g6574);
  not NOT_3181(g11237,II18163);
  not NOT_3182(II18166,g5778);
  not NOT_3183(g11240,II18166);
  not NOT_3184(II18169,g7195);
  not NOT_3185(g11243,II18169);
  not NOT_3186(II18172,g3722);
  not NOT_3187(g11246,II18172);
  not NOT_3188(II18175,g7085);
  not NOT_3189(g11249,II18175);
  not NOT_3190(II18178,g6838);
  not NOT_3191(g11252,II18178);
  not NOT_3192(II18181,g5636);
  not NOT_3193(g11255,II18181);
  not NOT_3194(II18184,g5837);
  not NOT_3195(g11256,II18184);
  not NOT_3196(II18187,g7391);
  not NOT_3197(g11259,II18187);
  not NOT_3198(II18211,g6232);
  not NOT_3199(g11265,II18211);
  not NOT_3200(II18214,g3254);
  not NOT_3201(g11268,II18214);
  not NOT_3202(II18217,g6314);
  not NOT_3203(g11271,II18217);
  not NOT_3204(II18220,g6232);
  not NOT_3205(g11274,II18220);
  not NOT_3206(II18223,g6448);
  not NOT_3207(g11277,II18223);
  not NOT_3208(II18226,g5668);
  not NOT_3209(g11278,II18226);
  not NOT_3210(II18229,g3410);
  not NOT_3211(g11281,II18229);
  not NOT_3212(II18232,g6519);
  not NOT_3213(g11284,II18232);
  not NOT_3214(II18235,g6369);
  not NOT_3215(g11287,II18235);
  not NOT_3216(II18238,g5593);
  not NOT_3217(g11290,II18238);
  not NOT_3218(II18241,g6713);
  not NOT_3219(g11291,II18241);
  not NOT_3220(II18244,g5720);
  not NOT_3221(g11294,II18244);
  not NOT_3222(II18247,g6945);
  not NOT_3223(g11297,II18247);
  not NOT_3224(II18250,g3566);
  not NOT_3225(g11300,II18250);
  not NOT_3226(II18253,g6783);
  not NOT_3227(g11303,II18253);
  not NOT_3228(II18256,g6574);
  not NOT_3229(g11306,II18256);
  not NOT_3230(II18259,g5778);
  not NOT_3231(g11309,II18259);
  not NOT_3232(II18262,g7195);
  not NOT_3233(g11312,II18262);
  not NOT_3234(II18265,g3722);
  not NOT_3235(g11315,II18265);
  not NOT_3236(II18268,g7085);
  not NOT_3237(g11318,II18268);
  not NOT_3238(II18271,g6838);
  not NOT_3239(g11321,II18271);
  not NOT_3240(II18274,g5837);
  not NOT_3241(g11324,II18274);
  not NOT_3242(II18277,g7391);
  not NOT_3243(g11327,II18277);
  not NOT_3244(g11332,g4094);
  not NOT_3245(II18295,g6314);
  not NOT_3246(g11341,II18295);
  not NOT_3247(II18298,g6232);
  not NOT_3248(g11344,II18298);
  not NOT_3249(II18302,g3254);
  not NOT_3250(g11348,II18302);
  not NOT_3251(II18305,g6314);
  not NOT_3252(g11351,II18305);
  not NOT_3253(II18308,g6448);
  not NOT_3254(g11354,II18308);
  not NOT_3255(II18311,g5668);
  not NOT_3256(g11355,II18311);
  not NOT_3257(II18314,g6369);
  not NOT_3258(g11358,II18314);
  not NOT_3259(II18317,g3410);
  not NOT_3260(g11361,II18317);
  not NOT_3261(II18320,g6519);
  not NOT_3262(g11364,II18320);
  not NOT_3263(II18323,g6369);
  not NOT_3264(g11367,II18323);
  not NOT_3265(II18326,g6713);
  not NOT_3266(g11370,II18326);
  not NOT_3267(II18329,g5720);
  not NOT_3268(g11373,II18329);
  not NOT_3269(II18332,g3566);
  not NOT_3270(g11376,II18332);
  not NOT_3271(II18335,g6783);
  not NOT_3272(g11379,II18335);
  not NOT_3273(II18338,g6574);
  not NOT_3274(g11382,II18338);
  not NOT_3275(II18341,g5610);
  not NOT_3276(g11385,II18341);
  not NOT_3277(II18344,g7015);
  not NOT_3278(g11386,II18344);
  not NOT_3279(II18347,g5778);
  not NOT_3280(g11389,II18347);
  not NOT_3281(II18350,g7195);
  not NOT_3282(g11392,II18350);
  not NOT_3283(II18353,g3722);
  not NOT_3284(g11395,II18353);
  not NOT_3285(II18356,g7085);
  not NOT_3286(g11398,II18356);
  not NOT_3287(II18359,g6838);
  not NOT_3288(g11401,II18359);
  not NOT_3289(II18362,g5837);
  not NOT_3290(g11404,II18362);
  not NOT_3291(II18365,g7391);
  not NOT_3292(g11407,II18365);
  not NOT_3293(II18375,g3254);
  not NOT_3294(g11411,II18375);
  not NOT_3295(II18378,g6314);
  not NOT_3296(g11414,II18378);
  not NOT_3297(II18381,g6232);
  not NOT_3298(g11417,II18381);
  not NOT_3299(II18386,g3254);
  not NOT_3300(g11422,II18386);
  not NOT_3301(II18389,g6519);
  not NOT_3302(g11425,II18389);
  not NOT_3303(II18392,g6369);
  not NOT_3304(g11428,II18392);
  not NOT_3305(II18396,g3410);
  not NOT_3306(g11432,II18396);
  not NOT_3307(II18399,g6519);
  not NOT_3308(g11435,II18399);
  not NOT_3309(II18402,g6713);
  not NOT_3310(g11438,II18402);
  not NOT_3311(II18405,g5720);
  not NOT_3312(g11441,II18405);
  not NOT_3313(II18408,g6574);
  not NOT_3314(g11444,II18408);
  not NOT_3315(II18411,g3566);
  not NOT_3316(g11447,II18411);
  not NOT_3317(II18414,g6783);
  not NOT_3318(g11450,II18414);
  not NOT_3319(II18417,g6574);
  not NOT_3320(g11453,II18417);
  not NOT_3321(II18420,g7015);
  not NOT_3322(g11456,II18420);
  not NOT_3323(II18423,g5778);
  not NOT_3324(g11459,II18423);
  not NOT_3325(II18426,g3722);
  not NOT_3326(g11462,II18426);
  not NOT_3327(II18429,g7085);
  not NOT_3328(g11465,II18429);
  not NOT_3329(II18432,g6838);
  not NOT_3330(g11468,II18432);
  not NOT_3331(II18435,g5635);
  not NOT_3332(g11471,II18435);
  not NOT_3333(II18438,g7265);
  not NOT_3334(g11472,II18438);
  not NOT_3335(II18441,g5837);
  not NOT_3336(g11475,II18441);
  not NOT_3337(II18444,g7391);
  not NOT_3338(g11478,II18444);
  not NOT_3339(g11481,g4204);
  not NOT_3340(g11490,g8276);
  not NOT_3341(II18449,g10868);
  not NOT_3342(g11491,II18449);
  not NOT_3343(II18452,g10930);
  not NOT_3344(g11492,II18452);
  not NOT_3345(II18455,g11031);
  not NOT_3346(g11493,II18455);
  not NOT_3347(II18458,g11208);
  not NOT_3348(g11494,II18458);
  not NOT_3349(II18461,g10931);
  not NOT_3350(g11495,II18461);
  not NOT_3351(II18464,g8620);
  not NOT_3352(g11496,II18464);
  not NOT_3353(II18467,g8769);
  not NOT_3354(g11497,II18467);
  not NOT_3355(II18470,g8808);
  not NOT_3356(g11498,II18470);
  not NOT_3357(II18473,g8839);
  not NOT_3358(g11499,II18473);
  not NOT_3359(II18476,g8791);
  not NOT_3360(g11500,II18476);
  not NOT_3361(II18479,g8820);
  not NOT_3362(g11501,II18479);
  not NOT_3363(II18482,g8859);
  not NOT_3364(g11502,II18482);
  not NOT_3365(II18485,g8809);
  not NOT_3366(g11503,II18485);
  not NOT_3367(II18488,g8840);
  not NOT_3368(g11504,II18488);
  not NOT_3369(II18491,g8891);
  not NOT_3370(g11505,II18491);
  not NOT_3371(II18494,g8821);
  not NOT_3372(g11506,II18494);
  not NOT_3373(II18497,g8860);
  not NOT_3374(g11507,II18497);
  not NOT_3375(II18500,g8924);
  not NOT_3376(g11508,II18500);
  not NOT_3377(II18503,g8658);
  not NOT_3378(g11509,II18503);
  not NOT_3379(II18506,g8699);
  not NOT_3380(g11510,II18506);
  not NOT_3381(II18509,g8770);
  not NOT_3382(g11511,II18509);
  not NOT_3383(II18512,g9309);
  not NOT_3384(g11512,II18512);
  not NOT_3385(II18515,g8843);
  not NOT_3386(g11513,II18515);
  not NOT_3387(II18518,g8893);
  not NOT_3388(g11514,II18518);
  not NOT_3389(II18521,g9449);
  not NOT_3390(g11515,II18521);
  not NOT_3391(II18524,g9640);
  not NOT_3392(g11516,II18524);
  not NOT_3393(II18527,g10017);
  not NOT_3394(g11517,II18527);
  not NOT_3395(II18530,g10888);
  not NOT_3396(g11518,II18530);
  not NOT_3397(II18533,g10967);
  not NOT_3398(g11519,II18533);
  not NOT_3399(II18536,g11101);
  not NOT_3400(g11520,II18536);
  not NOT_3401(II18539,g11290);
  not NOT_3402(g11521,II18539);
  not NOT_3403(II18542,g10968);
  not NOT_3404(g11522,II18542);
  not NOT_3405(II18545,g8630);
  not NOT_3406(g11523,II18545);
  not NOT_3407(II18548,g8792);
  not NOT_3408(g11524,II18548);
  not NOT_3409(II18551,g8824);
  not NOT_3410(g11525,II18551);
  not NOT_3411(II18554,g8866);
  not NOT_3412(g11526,II18554);
  not NOT_3413(II18557,g8810);
  not NOT_3414(g11527,II18557);
  not NOT_3415(II18560,g8844);
  not NOT_3416(g11528,II18560);
  not NOT_3417(II18563,g8897);
  not NOT_3418(g11529,II18563);
  not NOT_3419(II18566,g8825);
  not NOT_3420(g11530,II18566);
  not NOT_3421(II18569,g8867);
  not NOT_3422(g11531,II18569);
  not NOT_3423(II18572,g8931);
  not NOT_3424(g11532,II18572);
  not NOT_3425(II18575,g8845);
  not NOT_3426(g11533,II18575);
  not NOT_3427(II18578,g8898);
  not NOT_3428(g11534,II18578);
  not NOT_3429(II18581,g8964);
  not NOT_3430(g11535,II18581);
  not NOT_3431(II18584,g8677);
  not NOT_3432(g11536,II18584);
  not NOT_3433(II18587,g8718);
  not NOT_3434(g11537,II18587);
  not NOT_3435(II18590,g8793);
  not NOT_3436(g11538,II18590);
  not NOT_3437(II18593,g9390);
  not NOT_3438(g11539,II18593);
  not NOT_3439(II18596,g8870);
  not NOT_3440(g11540,II18596);
  not NOT_3441(II18599,g8933);
  not NOT_3442(g11541,II18599);
  not NOT_3443(II18602,g9591);
  not NOT_3444(g11542,II18602);
  not NOT_3445(II18605,g9786);
  not NOT_3446(g11543,II18605);
  not NOT_3447(II18608,g10126);
  not NOT_3448(g11544,II18608);
  not NOT_3449(II18611,g10909);
  not NOT_3450(g11545,II18611);
  not NOT_3451(II18614,g11002);
  not NOT_3452(g11546,II18614);
  not NOT_3453(II18617,g11169);
  not NOT_3454(g11547,II18617);
  not NOT_3455(II18620,g11385);
  not NOT_3456(g11548,II18620);
  not NOT_3457(II18623,g11003);
  not NOT_3458(g11549,II18623);
  not NOT_3459(II18626,g8649);
  not NOT_3460(g11550,II18626);
  not NOT_3461(II18629,g8811);
  not NOT_3462(g11551,II18629);
  not NOT_3463(II18632,g8850);
  not NOT_3464(g11552,II18632);
  not NOT_3465(II18635,g8904);
  not NOT_3466(g11553,II18635);
  not NOT_3467(II18638,g8826);
  not NOT_3468(g11554,II18638);
  not NOT_3469(II18641,g8871);
  not NOT_3470(g11555,II18641);
  not NOT_3471(II18644,g8937);
  not NOT_3472(g11556,II18644);
  not NOT_3473(II18647,g8851);
  not NOT_3474(g11557,II18647);
  not NOT_3475(II18650,g8905);
  not NOT_3476(g11558,II18650);
  not NOT_3477(II18653,g8971);
  not NOT_3478(g11559,II18653);
  not NOT_3479(II18656,g8872);
  not NOT_3480(g11560,II18656);
  not NOT_3481(II18659,g8938);
  not NOT_3482(g11561,II18659);
  not NOT_3483(II18662,g8996);
  not NOT_3484(g11562,II18662);
  not NOT_3485(II18665,g8689);
  not NOT_3486(g11563,II18665);
  not NOT_3487(II18668,g8756);
  not NOT_3488(g11564,II18668);
  not NOT_3489(II18671,g8812);
  not NOT_3490(g11565,II18671);
  not NOT_3491(II18674,g9487);
  not NOT_3492(g11566,II18674);
  not NOT_3493(II18677,g8908);
  not NOT_3494(g11567,II18677);
  not NOT_3495(II18680,g8973);
  not NOT_3496(g11568,II18680);
  not NOT_3497(II18683,g9733);
  not NOT_3498(g11569,II18683);
  not NOT_3499(II18686,g9932);
  not NOT_3500(g11570,II18686);
  not NOT_3501(II18689,g10231);
  not NOT_3502(g11571,II18689);
  not NOT_3503(II18692,g10935);
  not NOT_3504(g11572,II18692);
  not NOT_3505(II18695,g11054);
  not NOT_3506(g11573,II18695);
  not NOT_3507(II18698,g11255);
  not NOT_3508(g11574,II18698);
  not NOT_3509(II18701,g11471);
  not NOT_3510(g11575,II18701);
  not NOT_3511(II18704,g11055);
  not NOT_3512(g11576,II18704);
  not NOT_3513(II18707,g8665);
  not NOT_3514(g11577,II18707);
  not NOT_3515(II18710,g8827);
  not NOT_3516(g11578,II18710);
  not NOT_3517(II18713,g8877);
  not NOT_3518(g11579,II18713);
  not NOT_3519(II18716,g8944);
  not NOT_3520(g11580,II18716);
  not NOT_3521(II18719,g8852);
  not NOT_3522(g11581,II18719);
  not NOT_3523(II18722,g8909);
  not NOT_3524(g11582,II18722);
  not NOT_3525(II18725,g8977);
  not NOT_3526(g11583,II18725);
  not NOT_3527(II18728,g8878);
  not NOT_3528(g11584,II18728);
  not NOT_3529(II18731,g8945);
  not NOT_3530(g11585,II18731);
  not NOT_3531(II18734,g9003);
  not NOT_3532(g11586,II18734);
  not NOT_3533(II18737,g8910);
  not NOT_3534(g11587,II18737);
  not NOT_3535(II18740,g8978);
  not NOT_3536(g11588,II18740);
  not NOT_3537(II18743,g9025);
  not NOT_3538(g11589,II18743);
  not NOT_3539(II18746,g8707);
  not NOT_3540(g11590,II18746);
  not NOT_3541(II18749,g8779);
  not NOT_3542(g11591,II18749);
  not NOT_3543(II18752,g8828);
  not NOT_3544(g11592,II18752);
  not NOT_3545(II18755,g9629);
  not NOT_3546(g11593,II18755);
  not NOT_3547(II18758,g8948);
  not NOT_3548(g11594,II18758);
  not NOT_3549(II18761,g9005);
  not NOT_3550(g11595,II18761);
  not NOT_3551(II18764,g9879);
  not NOT_3552(g11596,II18764);
  not NOT_3553(II18767,g10086);
  not NOT_3554(g11597,II18767);
  not NOT_3555(II18770,g10333);
  not NOT_3556(g11598,II18770);
  not NOT_3557(II18773,g10830);
  not NOT_3558(g11599,II18773);
  not NOT_3559(II18777,g9050);
  not NOT_3560(g11603,II18777);
  not NOT_3561(II18780,g10870);
  not NOT_3562(g11606,II18780);
  not NOT_3563(II18784,g9067);
  not NOT_3564(g11608,II18784);
  not NOT_3565(II18787,g10910);
  not NOT_3566(g11611,II18787);
  not NOT_3567(II18791,g9084);
  not NOT_3568(g11613,II18791);
  not NOT_3569(II18794,g10973);
  not NOT_3570(g11616,II18794);
  not NOT_3571(g11620,g10601);
  not NOT_3572(g11623,g10961);
  not NOT_3573(II18810,g10813);
  not NOT_3574(g11628,II18810);
  not NOT_3575(II18813,g10850);
  not NOT_3576(g11629,II18813);
  not NOT_3577(II18817,g9067);
  not NOT_3578(g11633,II18817);
  not NOT_3579(II18820,g10890);
  not NOT_3580(g11636,II18820);
  not NOT_3581(II18824,g9084);
  not NOT_3582(g11638,II18824);
  not NOT_3583(II18827,g10936);
  not NOT_3584(g11641,II18827);
  not NOT_3585(g11642,g10646);
  not NOT_3586(II18835,g10834);
  not NOT_3587(g11651,II18835);
  not NOT_3588(II18838,g10871);
  not NOT_3589(g11652,II18838);
  not NOT_3590(II18842,g9084);
  not NOT_3591(g11656,II18842);
  not NOT_3592(II18845,g10911);
  not NOT_3593(g11659,II18845);
  not NOT_3594(II18854,g10854);
  not NOT_3595(g11670,II18854);
  not NOT_3596(II18857,g10891);
  not NOT_3597(g11671,II18857);
  not NOT_3598(II18866,g10875);
  not NOT_3599(g11682,II18866);
  not NOT_3600(g11706,g10928);
  not NOT_3601(g11732,g10826);
  not NOT_3602(g11734,g10843);
  not NOT_3603(g11735,g10859);
  not NOT_3604(g11736,g10862);
  not NOT_3605(g11737,g10809);
  not NOT_3606(g11740,g10877);
  not NOT_3607(g11741,g10880);
  not NOT_3608(g11742,g10883);
  not NOT_3609(g11743,g8530);
  not NOT_3610(g11745,g10892);
  not NOT_3611(g11746,g10895);
  not NOT_3612(g11747,g10898);
  not NOT_3613(g11748,g10901);
  not NOT_3614(II18929,g10711);
  not NOT_3615(g11749,II18929);
  not NOT_3616(g11758,g8514);
  not NOT_3617(g11761,g10912);
  not NOT_3618(g11762,g10915);
  not NOT_3619(g11763,g10918);
  not NOT_3620(g11764,g10921);
  not NOT_3621(g11765,g10924);
  not NOT_3622(g11766,g10886);
  not NOT_3623(II18943,g9149);
  not NOT_3624(g11769,II18943);
  not NOT_3625(g11770,g10932);
  not NOT_3626(g11774,g10937);
  not NOT_3627(g11775,g10940);
  not NOT_3628(g11776,g10943);
  not NOT_3629(g11777,g10946);
  not NOT_3630(g11778,g10949);
  not NOT_3631(g11779,g10906);
  not NOT_3632(g11782,g10963);
  not NOT_3633(g11783,g10966);
  not NOT_3634(II18962,g9159);
  not NOT_3635(g11786,II18962);
  not NOT_3636(g11787,g10969);
  not NOT_3637(II18969,g8726);
  not NOT_3638(g11791,II18969);
  not NOT_3639(g11794,g10974);
  not NOT_3640(g11795,g10977);
  not NOT_3641(g11796,g10980);
  not NOT_3642(g11797,g10983);
  not NOT_3643(g11798,g10867);
  not NOT_3644(g11801,g10988);
  not NOT_3645(g11802,g10991);
  not NOT_3646(g11803,g10994);
  not NOT_3647(g11804,g10995);
  not NOT_3648(g11808,g10996);
  not NOT_3649(g11809,g10999);
  not NOT_3650(II18990,g9183);
  not NOT_3651(g11812,II18990);
  not NOT_3652(g11813,g11004);
  not NOT_3653(g11817,g11008);
  not NOT_3654(g11818,g11011);
  not NOT_3655(g11819,g11014);
  not NOT_3656(g11820,g11017);
  not NOT_3657(g11821,g10848);
  not NOT_3658(g11824,g11022);
  not NOT_3659(g11825,g11025);
  not NOT_3660(g11826,g11028);
  not NOT_3661(g11827,g11032);
  not NOT_3662(g11829,g11035);
  not NOT_3663(g11834,g11036);
  not NOT_3664(g11835,g11039);
  not NOT_3665(g11836,g11042);
  not NOT_3666(g11837,g11045);
  not NOT_3667(g11841,g11048);
  not NOT_3668(g11842,g11051);
  not NOT_3669(II19025,g9225);
  not NOT_3670(g11845,II19025);
  not NOT_3671(g11846,g11056);
  not NOT_3672(II19030,g8726);
  not NOT_3673(g11848,II19030);
  not NOT_3674(g11852,g11063);
  not NOT_3675(g11853,g11066);
  not NOT_3676(g11854,g11078);
  not NOT_3677(g11856,g11079);
  not NOT_3678(g11857,g11082);
  not NOT_3679(g11858,g11085);
  not NOT_3680(g11859,g11088);
  not NOT_3681(g11862,g11091);
  not NOT_3682(g11866,g11092);
  not NOT_3683(g11867,g11095);
  not NOT_3684(g11868,g11098);
  not NOT_3685(g11869,g11102);
  not NOT_3686(g11871,g11105);
  not NOT_3687(g11876,g11108);
  not NOT_3688(g11877,g11111);
  not NOT_3689(g11878,g11114);
  not NOT_3690(g11879,g11117);
  not NOT_3691(g11883,g11120);
  not NOT_3692(g11884,g11123);
  not NOT_3693(g11886,g11126);
  not NOT_3694(g11887,g11129);
  not NOT_3695(g11888,g11021);
  not NOT_3696(g11891,g11132);
  not NOT_3697(g11892,g11135);
  not NOT_3698(g11893,g11138);
  not NOT_3699(g11894,g11141);
  not NOT_3700(g11895,g11144);
  not NOT_3701(g11898,g11145);
  not NOT_3702(g11899,g11148);
  not NOT_3703(g11900,g11151);
  not NOT_3704(g11901,g11154);
  not NOT_3705(g11904,g11157);
  not NOT_3706(g11908,g11160);
  not NOT_3707(g11909,g11163);
  not NOT_3708(g11910,g11166);
  not NOT_3709(g11911,g11170);
  not NOT_3710(g11913,g11173);
  not NOT_3711(g11918,g11176);
  not NOT_3712(g11919,g11179);
  not NOT_3713(g11920,g11182);
  not NOT_3714(g11921,g11185);
  not NOT_3715(II19105,g8726);
  not NOT_3716(g11923,II19105);
  not NOT_3717(g11927,g10987);
  not NOT_3718(g11929,g11199);
  not NOT_3719(g11930,g11202);
  not NOT_3720(g11931,g11205);
  not NOT_3721(g11932,g11209);
  not NOT_3722(g11933,g11210);
  not NOT_3723(g11936,g11213);
  not NOT_3724(II19119,g9202);
  not NOT_3725(g11937,II19119);
  not NOT_3726(g11941,g11216);
  not NOT_3727(g11942,g11219);
  not NOT_3728(g11943,g11222);
  not NOT_3729(g11944,g11225);
  not NOT_3730(g11945,g11228);
  not NOT_3731(g11948,g11231);
  not NOT_3732(g11949,g11234);
  not NOT_3733(g11950,g11237);
  not NOT_3734(g11951,g11240);
  not NOT_3735(g11954,g11243);
  not NOT_3736(g11958,g11246);
  not NOT_3737(g11959,g11249);
  not NOT_3738(g11960,g11252);
  not NOT_3739(g11961,g11256);
  not NOT_3740(g11963,g11259);
  not NOT_3741(g11968,g11265);
  not NOT_3742(g11969,g11268);
  not NOT_3743(g11970,g11271);
  not NOT_3744(g11971,g11274);
  not NOT_3745(g11972,g11277);
  not NOT_3746(g11973,g11278);
  not NOT_3747(II19160,g10549);
  not NOT_3748(g11976,II19160);
  not NOT_3749(g11982,g11281);
  not NOT_3750(g11983,g11284);
  not NOT_3751(g11984,g11287);
  not NOT_3752(g11985,g11291);
  not NOT_3753(g11986,g11294);
  not NOT_3754(g11989,g11297);
  not NOT_3755(II19174,g9263);
  not NOT_3756(g11990,II19174);
  not NOT_3757(g11994,g11300);
  not NOT_3758(g11995,g11303);
  not NOT_3759(g11996,g11306);
  not NOT_3760(g11997,g11309);
  not NOT_3761(g11998,g11312);
  not NOT_3762(g12001,g11315);
  not NOT_3763(g12002,g11318);
  not NOT_3764(g12003,g11321);
  not NOT_3765(g12004,g11324);
  not NOT_3766(g12007,g11327);
  not NOT_3767(II19195,g8726);
  not NOT_3768(g12009,II19195);
  not NOT_3769(g12013,g10772);
  not NOT_3770(g12017,g10100);
  not NOT_3771(g12020,g11341);
  not NOT_3772(g12021,g11344);
  not NOT_3773(g12022,g11348);
  not NOT_3774(g12023,g11351);
  not NOT_3775(g12024,g11354);
  not NOT_3776(g12025,g11355);
  not NOT_3777(II19208,g10424);
  not NOT_3778(g12027,II19208);
  not NOT_3779(II19211,g10486);
  not NOT_3780(g12030,II19211);
  not NOT_3781(g12037,g11358);
  not NOT_3782(g12038,g11361);
  not NOT_3783(g12039,g11364);
  not NOT_3784(g12040,g11367);
  not NOT_3785(g12041,g11370);
  not NOT_3786(g12042,g11373);
  not NOT_3787(II19226,g10606);
  not NOT_3788(g12045,II19226);
  not NOT_3789(g12051,g11376);
  not NOT_3790(g12052,g11379);
  not NOT_3791(g12053,g11382);
  not NOT_3792(g12054,g11386);
  not NOT_3793(g12055,g11389);
  not NOT_3794(g12058,g11392);
  not NOT_3795(II19240,g9341);
  not NOT_3796(g12059,II19240);
  not NOT_3797(g12063,g11395);
  not NOT_3798(g12064,g11398);
  not NOT_3799(g12065,g11401);
  not NOT_3800(g12066,g11404);
  not NOT_3801(g12067,g11407);
  not NOT_3802(g12071,g10783);
  not NOT_3803(g12075,g11411);
  not NOT_3804(g12076,g11414);
  not NOT_3805(g12077,g11417);
  not NOT_3806(g12078,g11422);
  not NOT_3807(g12084,g11425);
  not NOT_3808(g12085,g11428);
  not NOT_3809(g12086,g11432);
  not NOT_3810(g12087,g11435);
  not NOT_3811(g12088,g11438);
  not NOT_3812(g12089,g11441);
  not NOT_3813(II19271,g10500);
  not NOT_3814(g12091,II19271);
  not NOT_3815(II19274,g10560);
  not NOT_3816(g12094,II19274);
  not NOT_3817(g12101,g11444);
  not NOT_3818(g12102,g11447);
  not NOT_3819(g12103,g11450);
  not NOT_3820(g12104,g11453);
  not NOT_3821(g12105,g11456);
  not NOT_3822(g12106,g11459);
  not NOT_3823(II19289,g10653);
  not NOT_3824(g12109,II19289);
  not NOT_3825(g12115,g11462);
  not NOT_3826(g12116,g11465);
  not NOT_3827(g12117,g11468);
  not NOT_3828(g12118,g11472);
  not NOT_3829(g12119,g11475);
  not NOT_3830(g12122,g11478);
  not NOT_3831(II19303,g9422);
  not NOT_3832(g12123,II19303);
  not NOT_3833(II19307,g8726);
  not NOT_3834(g12125,II19307);
  not NOT_3835(g12130,g10788);
  not NOT_3836(g12134,g8321);
  not NOT_3837(g12135,g8324);
  not NOT_3838(II19315,g10424);
  not NOT_3839(g12136,II19315);
  not NOT_3840(II19318,g10486);
  not NOT_3841(g12139,II19318);
  not NOT_3842(II19321,g10549);
  not NOT_3843(g12142,II19321);
  not NOT_3844(g12147,g8330);
  not NOT_3845(g12148,g8333);
  not NOT_3846(g12149,g8336);
  not NOT_3847(g12150,g8341);
  not NOT_3848(g12156,g8344);
  not NOT_3849(g12157,g8347);
  not NOT_3850(g12158,g8351);
  not NOT_3851(g12159,g8354);
  not NOT_3852(g12160,g8357);
  not NOT_3853(g12161,g8360);
  not NOT_3854(II19342,g10574);
  not NOT_3855(g12163,II19342);
  not NOT_3856(II19345,g10617);
  not NOT_3857(g12166,II19345);
  not NOT_3858(g12173,g8363);
  not NOT_3859(g12174,g8366);
  not NOT_3860(g12175,g8369);
  not NOT_3861(g12176,g8372);
  not NOT_3862(g12177,g8375);
  not NOT_3863(g12178,g8378);
  not NOT_3864(II19360,g10683);
  not NOT_3865(g12181,II19360);
  not NOT_3866(g12187,g8285);
  not NOT_3867(g12191,g8382);
  not NOT_3868(g12196,g8388);
  not NOT_3869(g12197,g8391);
  not NOT_3870(II19374,g10500);
  not NOT_3871(g12198,II19374);
  not NOT_3872(II19377,g10560);
  not NOT_3873(g12201,II19377);
  not NOT_3874(II19380,g10606);
  not NOT_3875(g12204,II19380);
  not NOT_3876(g12209,g8397);
  not NOT_3877(g12210,g8400);
  not NOT_3878(g12211,g8403);
  not NOT_3879(g12212,g8408);
  not NOT_3880(g12218,g8411);
  not NOT_3881(g12219,g8414);
  not NOT_3882(g12220,g8418);
  not NOT_3883(g12221,g8421);
  not NOT_3884(g12222,g8424);
  not NOT_3885(g12223,g8427);
  not NOT_3886(II19401,g10631);
  not NOT_3887(g12225,II19401);
  not NOT_3888(II19404,g10664);
  not NOT_3889(g12228,II19404);
  not NOT_3890(g12235,g8294);
  not NOT_3891(II19412,g10486);
  not NOT_3892(g12239,II19412);
  not NOT_3893(II19415,g10549);
  not NOT_3894(g12242,II19415);
  not NOT_3895(g12246,g8434);
  not NOT_3896(g12251,g8440);
  not NOT_3897(g12252,g8443);
  not NOT_3898(II19426,g10574);
  not NOT_3899(g12253,II19426);
  not NOT_3900(II19429,g10617);
  not NOT_3901(g12256,II19429);
  not NOT_3902(II19432,g10653);
  not NOT_3903(g12259,II19432);
  not NOT_3904(g12264,g8449);
  not NOT_3905(g12265,g8452);
  not NOT_3906(g12266,g8455);
  not NOT_3907(g12267,g8460);
  not NOT_3908(g12275,g8303);
  not NOT_3909(II19449,g10424);
  not NOT_3910(g12279,II19449);
  not NOT_3911(II19452,g10560);
  not NOT_3912(g12282,II19452);
  not NOT_3913(II19455,g10606);
  not NOT_3914(g12285,II19455);
  not NOT_3915(g12289,g8469);
  not NOT_3916(g12294,g8475);
  not NOT_3917(g12295,g8478);
  not NOT_3918(II19466,g10631);
  not NOT_3919(g12296,II19466);
  not NOT_3920(II19469,g10664);
  not NOT_3921(g12299,II19469);
  not NOT_3922(II19472,g10683);
  not NOT_3923(g12302,II19472);
  not NOT_3924(g12308,g8312);
  not NOT_3925(II19479,g10549);
  not NOT_3926(g12312,II19479);
  not NOT_3927(II19482,g10500);
  not NOT_3928(g12315,II19482);
  not NOT_3929(II19485,g10617);
  not NOT_3930(g12318,II19485);
  not NOT_3931(II19488,g10653);
  not NOT_3932(g12321,II19488);
  not NOT_3933(g12325,g8494);
  not NOT_3934(g12332,g10829);
  not NOT_3935(II19500,g10424);
  not NOT_3936(g12333,II19500);
  not NOT_3937(II19503,g10486);
  not NOT_3938(g12336,II19503);
  not NOT_3939(II19507,g10606);
  not NOT_3940(g12340,II19507);
  not NOT_3941(II19510,g10574);
  not NOT_3942(g12343,II19510);
  not NOT_3943(II19513,g10664);
  not NOT_3944(g12346,II19513);
  not NOT_3945(II19516,g10683);
  not NOT_3946(g12349,II19516);
  not NOT_3947(g12354,g8381);
  not NOT_3948(g12362,g10866);
  not NOT_3949(II19523,g10500);
  not NOT_3950(g12363,II19523);
  not NOT_3951(II19526,g10560);
  not NOT_3952(g12366,II19526);
  not NOT_3953(II19530,g10653);
  not NOT_3954(g12370,II19530);
  not NOT_3955(II19533,g10631);
  not NOT_3956(g12373,II19533);
  not NOT_3957(g12378,g10847);
  not NOT_3958(II19539,g10549);
  not NOT_3959(g12379,II19539);
  not NOT_3960(II19542,g10574);
  not NOT_3961(g12382,II19542);
  not NOT_3962(II19545,g10617);
  not NOT_3963(g12385,II19545);
  not NOT_3964(II19549,g10683);
  not NOT_3965(g12389,II19549);
  not NOT_3966(II19552,g8430);
  not NOT_3967(g12392,II19552);
  not NOT_3968(g12408,g11020);
  not NOT_3969(II19557,g10606);
  not NOT_3970(g12409,II19557);
  not NOT_3971(II19560,g10631);
  not NOT_3972(g12412,II19560);
  not NOT_3973(II19563,g10664);
  not NOT_3974(g12415,II19563);
  not NOT_3975(g12420,g10986);
  not NOT_3976(II19569,g10653);
  not NOT_3977(g12421,II19569);
  not NOT_3978(g12424,g10962);
  not NOT_3979(II19573,g8835);
  not NOT_3980(g12425,II19573);
  not NOT_3981(II19576,g10683);
  not NOT_3982(g12426,II19576);
  not NOT_3983(g12430,g10905);
  not NOT_3984(II19582,g8862);
  not NOT_3985(g12432,II19582);
  not NOT_3986(g12434,g10929);
  not NOT_3987(II19587,g9173);
  not NOT_3988(g12435,II19587);
  not NOT_3989(II19591,g8900);
  not NOT_3990(g12437,II19591);
  not NOT_3991(g12438,g10846);
  not NOT_3992(II19595,g10810);
  not NOT_3993(g12439,II19595);
  not NOT_3994(II19598,g9215);
  not NOT_3995(g12440,II19598);
  not NOT_3996(II19602,g8940);
  not NOT_3997(g12442,II19602);
  not NOT_3998(II19605,g10797);
  not NOT_3999(g12443,II19605);
  not NOT_4000(II19608,g10831);
  not NOT_4001(g12444,II19608);
  not NOT_4002(II19611,g9276);
  not NOT_4003(g12445,II19611);
  not NOT_4004(II19615,g10789);
  not NOT_4005(g12447,II19615);
  not NOT_4006(II19618,g10814);
  not NOT_4007(g12448,II19618);
  not NOT_4008(II19621,g10851);
  not NOT_4009(g12449,II19621);
  not NOT_4010(II19624,g9354);
  not NOT_4011(g12450,II19624);
  not NOT_4012(II19628,g10784);
  not NOT_4013(g12452,II19628);
  not NOT_4014(II19631,g10801);
  not NOT_4015(g12453,II19631);
  not NOT_4016(II19634,g10835);
  not NOT_4017(g12454,II19634);
  not NOT_4018(II19637,g10872);
  not NOT_4019(g12455,II19637);
  not NOT_4020(g12456,g8602);
  not NOT_4021(II19642,g10793);
  not NOT_4022(g12460,II19642);
  not NOT_4023(II19645,g10818);
  not NOT_4024(g12461,II19645);
  not NOT_4025(II19648,g10855);
  not NOT_4026(g12462,II19648);
  not NOT_4027(g12463,g10730);
  not NOT_4028(g12466,g8614);
  not NOT_4029(II19654,g10805);
  not NOT_4030(g12470,II19654);
  not NOT_4031(II19657,g10839);
  not NOT_4032(g12471,II19657);
  not NOT_4033(g12472,g8617);
  not NOT_4034(g12473,g8580);
  not NOT_4035(g12476,g8622);
  not NOT_4036(g12478,g10749);
  not NOT_4037(g12481,g8627);
  not NOT_4038(II19667,g10822);
  not NOT_4039(g12485,II19667);
  not NOT_4040(g12490,g8587);
  not NOT_4041(g12493,g8632);
  not NOT_4042(g12495,g10767);
  not NOT_4043(g12498,g8637);
  not NOT_4044(g12502,g8640);
  not NOT_4045(g12504,g8643);
  not NOT_4046(g12505,g8646);
  not NOT_4047(g12510,g8594);
  not NOT_4048(g12513,g8651);
  not NOT_4049(g12515,g10773);
  not NOT_4050(g12518,g8655);
  not NOT_4051(II19689,g10016);
  not NOT_4052(g12519,II19689);
  not NOT_4053(g12521,g8659);
  not NOT_4054(g12522,g8662);
  not NOT_4055(g12527,g8605);
  not NOT_4056(g12530,g8667);
  not NOT_4057(g12532,g8670);
  not NOT_4058(g12533,g8673);
  not NOT_4059(II19702,g10125);
  not NOT_4060(g12534,II19702);
  not NOT_4061(g12536,g8678);
  not NOT_4062(g12537,g8681);
  not NOT_4063(g12542,g8684);
  not NOT_4064(II19711,g10230);
  not NOT_4065(g12543,II19711);
  not NOT_4066(g12545,g8690);
  not NOT_4067(g12546,g8693);
  not NOT_4068(g12547,g8696);
  not NOT_4069(II19718,g8726);
  not NOT_4070(g12548,II19718);
  not NOT_4071(g12551,g8700);
  not NOT_4072(II19722,g10332);
  not NOT_4073(g12552,II19722);
  not NOT_4074(g12553,g8708);
  not NOT_4075(g12554,g8711);
  not NOT_4076(II19727,g8726);
  not NOT_4077(g12555,II19727);
  not NOT_4078(g12558,g8714);
  not NOT_4079(g12559,g8719);
  not NOT_4080(g12560,g8745);
  not NOT_4081(II19733,g8726);
  not NOT_4082(g12561,II19733);
  not NOT_4083(II19736,g9184);
  not NOT_4084(g12564,II19736);
  not NOT_4085(II19739,g10694);
  not NOT_4086(g12565,II19739);
  not NOT_4087(g12596,g8748);
  not NOT_4088(g12597,g8752);
  not NOT_4089(g12598,g8757);
  not NOT_4090(g12599,g8763);
  not NOT_4091(g12600,g8766);
  not NOT_4092(II19747,g8726);
  not NOT_4093(g12601,II19747);
  not NOT_4094(II19750,g8726);
  not NOT_4095(g12604,II19750);
  not NOT_4096(II19753,g9229);
  not NOT_4097(g12607,II19753);
  not NOT_4098(II19756,g10424);
  not NOT_4099(g12608,II19756);
  not NOT_4100(II19759,g10714);
  not NOT_4101(g12611,II19759);
  not NOT_4102(g12642,g8771);
  not NOT_4103(g12643,g8775);
  not NOT_4104(g12644,g8780);
  not NOT_4105(g12645,g8785);
  not NOT_4106(g12646,g8788);
  not NOT_4107(II19767,g8726);
  not NOT_4108(g12647,II19767);
  not NOT_4109(II19771,g10038);
  not NOT_4110(g12651,II19771);
  not NOT_4111(II19774,g10500);
  not NOT_4112(g12654,II19774);
  not NOT_4113(II19777,g10735);
  not NOT_4114(g12657,II19777);
  not NOT_4115(g12688,g8794);
  not NOT_4116(g12689,g8798);
  not NOT_4117(g12690,g8802);
  not NOT_4118(g12691,g8805);
  not NOT_4119(II19784,g8726);
  not NOT_4120(g12692,II19784);
  not NOT_4121(II19787,g8726);
  not NOT_4122(g12695,II19787);
  not NOT_4123(II19791,g10486);
  not NOT_4124(g12699,II19791);
  not NOT_4125(II19794,g10676);
  not NOT_4126(g12702,II19794);
  not NOT_4127(II19797,g10147);
  not NOT_4128(g12705,II19797);
  not NOT_4129(II19800,g10574);
  not NOT_4130(g12708,II19800);
  not NOT_4131(II19803,g10754);
  not NOT_4132(g12711,II19803);
  not NOT_4133(g12742,g8813);
  not NOT_4134(g12743,g8817);
  not NOT_4135(II19808,g8726);
  not NOT_4136(g12744,II19808);
  not NOT_4137(g12748,g8823);
  not NOT_4138(II19813,g10649);
  not NOT_4139(g12749,II19813);
  not NOT_4140(II19816,g10703);
  not NOT_4141(g12752,II19816);
  not NOT_4142(II19820,g10560);
  not NOT_4143(g12756,II19820);
  not NOT_4144(II19823,g10705);
  not NOT_4145(g12759,II19823);
  not NOT_4146(II19826,g10252);
  not NOT_4147(g12762,II19826);
  not NOT_4148(II19829,g10631);
  not NOT_4149(g12765,II19829);
  not NOT_4150(g12768,g8829);
  not NOT_4151(II19833,g8726);
  not NOT_4152(g12769,II19833);
  not NOT_4153(II19836,g8726);
  not NOT_4154(g12772,II19836);
  not NOT_4155(g12775,g8832);
  not NOT_4156(g12776,g10766);
  not NOT_4157(g12782,g8836);
  not NOT_4158(II19844,g8533);
  not NOT_4159(g12783,II19844);
  not NOT_4160(II19847,g10677);
  not NOT_4161(g12786,II19847);
  not NOT_4162(g12790,g8847);
  not NOT_4163(II19852,g10679);
  not NOT_4164(g12791,II19852);
  not NOT_4165(II19855,g10723);
  not NOT_4166(g12794,II19855);
  not NOT_4167(II19859,g10617);
  not NOT_4168(g12798,II19859);
  not NOT_4169(II19862,g10725);
  not NOT_4170(g12801,II19862);
  not NOT_4171(II19865,g10354);
  not NOT_4172(g12804,II19865);
  not NOT_4173(g12807,g8853);
  not NOT_4174(II19869,g8726);
  not NOT_4175(g12808,II19869);
  not NOT_4176(II19872,g8317);
  not NOT_4177(g12811,II19872);
  not NOT_4178(g12815,g8856);
  not NOT_4179(II19877,g8547);
  not NOT_4180(g12816,II19877);
  not NOT_4181(g12821,g8863);
  not NOT_4182(II19883,g8550);
  not NOT_4183(g12822,II19883);
  not NOT_4184(II19886,g10706);
  not NOT_4185(g12825,II19886);
  not NOT_4186(g12829,g8874);
  not NOT_4187(II19891,g10708);
  not NOT_4188(g12830,II19891);
  not NOT_4189(II19894,g10744);
  not NOT_4190(g12833,II19894);
  not NOT_4191(II19898,g10664);
  not NOT_4192(g12837,II19898);
  not NOT_4193(II19901,g10746);
  not NOT_4194(g12840,II19901);
  not NOT_4195(g12843,g8879);
  not NOT_4196(II19905,g8726);
  not NOT_4197(g12844,II19905);
  not NOT_4198(g12847,g8882);
  not NOT_4199(g12848,g11059);
  not NOT_4200(g12850,g8885);
  not NOT_4201(g12851,g8888);
  not NOT_4202(g12853,g8894);
  not NOT_4203(II19915,g8560);
  not NOT_4204(g12854,II19915);
  not NOT_4205(g12859,g8901);
  not NOT_4206(II19921,g8563);
  not NOT_4207(g12860,II19921);
  not NOT_4208(II19924,g10726);
  not NOT_4209(g12863,II19924);
  not NOT_4210(g12867,g8912);
  not NOT_4211(II19929,g10728);
  not NOT_4212(g12868,II19929);
  not NOT_4213(II19932,g10763);
  not NOT_4214(g12871,II19932);
  not NOT_4215(g12874,g8915);
  not NOT_4216(g12875,g10779);
  not NOT_4217(g12881,g8918);
  not NOT_4218(g12882,g8921);
  not NOT_4219(g12891,g8925);
  not NOT_4220(g12892,g8928);
  not NOT_4221(g12894,g8934);
  not NOT_4222(II19952,g8571);
  not NOT_4223(g12895,II19952);
  not NOT_4224(g12900,g8941);
  not NOT_4225(II19958,g8574);
  not NOT_4226(g12901,II19958);
  not NOT_4227(II19961,g10747);
  not NOT_4228(g12904,II19961);
  not NOT_4229(g12907,g8949);
  not NOT_4230(g12909,g10904);
  not NOT_4231(g12914,g8952);
  not NOT_4232(g12915,g8955);
  not NOT_4233(g12921,g8958);
  not NOT_4234(g12922,g8961);
  not NOT_4235(g12931,g8965);
  not NOT_4236(g12932,g8968);
  not NOT_4237(g12934,g8974);
  not NOT_4238(II19986,g8577);
  not NOT_4239(g12935,II19986);
  not NOT_4240(g12940,g8980);
  not NOT_4241(g12943,g8984);
  not NOT_4242(g12944,g8987);
  not NOT_4243(g12950,g8990);
  not NOT_4244(g12951,g8993);
  not NOT_4245(g12960,g8997);
  not NOT_4246(g12961,g9000);
  not NOT_4247(II20009,g8313);
  not NOT_4248(g12962,II20009);
  not NOT_4249(g12965,g9006);
  not NOT_4250(g12969,g9010);
  not NOT_4251(g12972,g9013);
  not NOT_4252(g12973,g9016);
  not NOT_4253(g12979,g9019);
  not NOT_4254(g12980,g9022);
  not NOT_4255(g12993,g9035);
  not NOT_4256(g12996,g9038);
  not NOT_4257(g12997,g9041);
  not NOT_4258(g12998,g9044);
  not NOT_4259(g13003,g9058);
  not NOT_4260(II20062,g10480);
  not NOT_4261(g13011,II20062);
  not NOT_4262(g13025,g10810);
  not NOT_4263(g13033,g10797);
  not NOT_4264(g13036,g10831);
  not NOT_4265(g13043,g10789);
  not NOT_4266(g13046,g10814);
  not NOT_4267(g13049,g10851);
  not NOT_4268(g13057,g10784);
  not NOT_4269(g13060,g10801);
  not NOT_4270(g13063,g10835);
  not NOT_4271(g13066,g10872);
  not NOT_4272(II20117,g10876);
  not NOT_4273(g13070,II20117);
  not NOT_4274(g13073,g10793);
  not NOT_4275(g13076,g10818);
  not NOT_4276(g13079,g10855);
  not NOT_4277(g13092,g10805);
  not NOT_4278(g13095,g10839);
  not NOT_4279(g13101,g9128);
  not NOT_4280(g13107,g10822);
  not NOT_4281(g13117,g9134);
  not NOT_4282(g13130,g9140);
  not NOT_4283(g13141,g9146);
  not NOT_4284(g13148,g9170);
  not NOT_4285(g13151,g9184);
  not NOT_4286(g13152,g9196);
  not NOT_4287(g13153,g9199);
  not NOT_4288(g13154,g9212);
  not NOT_4289(g13157,g9229);
  not NOT_4290(g13158,g9242);
  not NOT_4291(g13159,g9245);
  not NOT_4292(g13161,g9257);
  not NOT_4293(g13162,g9260);
  not NOT_4294(g13163,g9273);
  not NOT_4295(g13166,g9290);
  not NOT_4296(g13167,g9303);
  not NOT_4297(g13168,g9306);
  not NOT_4298(g13169,g9320);
  not NOT_4299(g13170,g9323);
  not NOT_4300(g13172,g9335);
  not NOT_4301(g13173,g9338);
  not NOT_4302(g13174,g9351);
  not NOT_4303(g13176,g9368);
  not NOT_4304(g13177,g9371);
  not NOT_4305(g13178,g9384);
  not NOT_4306(g13179,g9387);
  not NOT_4307(g13180,g9401);
  not NOT_4308(g13181,g9404);
  not NOT_4309(g13183,g9416);
  not NOT_4310(g13184,g9419);
  not NOT_4311(g13185,g9443);
  not NOT_4312(g13186,g9446);
  not NOT_4313(g13187,g9450);
  not NOT_4314(g13188,g9465);
  not NOT_4315(g13189,g9468);
  not NOT_4316(g13190,g9481);
  not NOT_4317(g13191,g9484);
  not NOT_4318(g13192,g9498);
  not NOT_4319(g13193,g9501);
  not NOT_4320(g13195,g9524);
  not NOT_4321(g13196,g9528);
  not NOT_4322(g13197,g9531);
  not NOT_4323(g13198,g9585);
  not NOT_4324(g13199,g9588);
  not NOT_4325(g13200,g9592);
  not NOT_4326(g13201,g9607);
  not NOT_4327(g13202,g9610);
  not NOT_4328(g13203,g9623);
  not NOT_4329(g13204,g9626);
  not NOT_4330(g13205,g9641);
  not NOT_4331(g13206,g9644);
  not NOT_4332(g13207,g9666);
  not NOT_4333(g13208,g9670);
  not NOT_4334(g13209,g9673);
  not NOT_4335(g13210,g9727);
  not NOT_4336(g13211,g9730);
  not NOT_4337(g13212,g9734);
  not NOT_4338(g13213,g9749);
  not NOT_4339(g13214,g9752);
  not NOT_4340(II20264,g9027);
  not NOT_4341(g13215,II20264);
  not NOT_4342(g13218,g9767);
  not NOT_4343(g13219,g9770);
  not NOT_4344(g13220,g9787);
  not NOT_4345(g13221,g9790);
  not NOT_4346(g13222,g9812);
  not NOT_4347(g13223,g9816);
  not NOT_4348(g13224,g9819);
  not NOT_4349(g13225,g9873);
  not NOT_4350(g13226,g9876);
  not NOT_4351(g13227,g9880);
  not NOT_4352(II20278,g9027);
  not NOT_4353(g13229,II20278);
  not NOT_4354(g13232,g9895);
  not NOT_4355(g13233,g9898);
  not NOT_4356(II20283,g9050);
  not NOT_4357(g13234,II20283);
  not NOT_4358(g13237,g9913);
  not NOT_4359(g13238,g9916);
  not NOT_4360(g13239,g9933);
  not NOT_4361(g13240,g9936);
  not NOT_4362(g13241,g9958);
  not NOT_4363(g13242,g9962);
  not NOT_4364(g13243,g9965);
  not NOT_4365(g13244,g10004);
  not NOT_4366(II20295,g10015);
  not NOT_4367(g13246,II20295);
  not NOT_4368(II20299,g10800);
  not NOT_4369(g13248,II20299);
  not NOT_4370(g13249,g10018);
  not NOT_4371(g13250,g10021);
  not NOT_4372(II20305,g9050);
  not NOT_4373(g13252,II20305);
  not NOT_4374(g13255,g10049);
  not NOT_4375(g13256,g10052);
  not NOT_4376(II20310,g9067);
  not NOT_4377(g13257,II20310);
  not NOT_4378(g13260,g10067);
  not NOT_4379(g13261,g10070);
  not NOT_4380(g13262,g10087);
  not NOT_4381(g13263,g10090);
  not NOT_4382(g13264,g10096);
  not NOT_4383(g13265,g8568);
  not NOT_4384(II20320,g10792);
  not NOT_4385(g13267,II20320);
  not NOT_4386(g13268,g10109);
  not NOT_4387(II20324,g10124);
  not NOT_4388(g13269,II20324);
  not NOT_4389(II20328,g10817);
  not NOT_4390(g13271,II20328);
  not NOT_4391(g13272,g10127);
  not NOT_4392(g13273,g10130);
  not NOT_4393(II20334,g9067);
  not NOT_4394(g13275,II20334);
  not NOT_4395(g13278,g10158);
  not NOT_4396(g13279,g10161);
  not NOT_4397(II20339,g9084);
  not NOT_4398(g13280,II20339);
  not NOT_4399(g13283,g10176);
  not NOT_4400(g13284,g10179);
  not NOT_4401(g13285,g10189);
  not NOT_4402(II20347,g10787);
  not NOT_4403(g13290,II20347);
  not NOT_4404(II20351,g10804);
  not NOT_4405(g13292,II20351);
  not NOT_4406(g13293,g10214);
  not NOT_4407(II20355,g10229);
  not NOT_4408(g13294,II20355);
  not NOT_4409(II20359,g10838);
  not NOT_4410(g13296,II20359);
  not NOT_4411(g13297,g10232);
  not NOT_4412(g13298,g10235);
  not NOT_4413(II20365,g9084);
  not NOT_4414(g13300,II20365);
  not NOT_4415(g13303,g10263);
  not NOT_4416(g13304,g10266);
  not NOT_4417(g13308,g10273);
  not NOT_4418(g13309,g10276);
  not NOT_4419(II20376,g8569);
  not NOT_4420(g13317,II20376);
  not NOT_4421(II20379,g11213);
  not NOT_4422(g13318,II20379);
  not NOT_4423(II20382,g10907);
  not NOT_4424(g13319,II20382);
  not NOT_4425(II20386,g10796);
  not NOT_4426(g13321,II20386);
  not NOT_4427(II20390,g10821);
  not NOT_4428(g13323,II20390);
  not NOT_4429(g13324,g10316);
  not NOT_4430(II20394,g10331);
  not NOT_4431(g13325,II20394);
  not NOT_4432(II20398,g10858);
  not NOT_4433(g13327,II20398);
  not NOT_4434(g13328,g10334);
  not NOT_4435(g13329,g10337);
  not NOT_4436(g13330,g10357);
  not NOT_4437(II20407,g9027);
  not NOT_4438(g13336,II20407);
  not NOT_4439(II20410,g10887);
  not NOT_4440(g13339,II20410);
  not NOT_4441(II20414,g8575);
  not NOT_4442(g13341,II20414);
  not NOT_4443(II20417,g10933);
  not NOT_4444(g13342,II20417);
  not NOT_4445(II20421,g10808);
  not NOT_4446(g13344,II20421);
  not NOT_4447(II20425,g10842);
  not NOT_4448(g13346,II20425);
  not NOT_4449(g13347,g10409);
  not NOT_4450(g13351,g10416);
  not NOT_4451(g13352,g10419);
  not NOT_4452(II20441,g9027);
  not NOT_4453(g13356,II20441);
  not NOT_4454(II20444,g10869);
  not NOT_4455(g13359,II20444);
  not NOT_4456(II20448,g9050);
  not NOT_4457(g13361,II20448);
  not NOT_4458(II20451,g10908);
  not NOT_4459(g13364,II20451);
  not NOT_4460(II20455,g8578);
  not NOT_4461(g13366,II20455);
  not NOT_4462(II20458,g10972);
  not NOT_4463(g13367,II20458);
  not NOT_4464(II20462,g10825);
  not NOT_4465(g13369,II20462);
  not NOT_4466(g13373,g10482);
  not NOT_4467(II20476,g9027);
  not NOT_4468(g13381,II20476);
  not NOT_4469(II20479,g10849);
  not NOT_4470(g13384,II20479);
  not NOT_4471(II20483,g9050);
  not NOT_4472(g13386,II20483);
  not NOT_4473(II20486,g10889);
  not NOT_4474(g13389,II20486);
  not NOT_4475(II20490,g9067);
  not NOT_4476(g13391,II20490);
  not NOT_4477(II20493,g10934);
  not NOT_4478(g13394,II20493);
  not NOT_4479(II20497,g8579);
  not NOT_4480(g13396,II20497);
  not NOT_4481(II20500,g11007);
  not NOT_4482(g13397,II20500);
  not NOT_4483(g13398,g10542);
  not NOT_4484(g13400,g10545);
  not NOT_4485(II20514,g11769);
  not NOT_4486(g13405,II20514);
  not NOT_4487(II20517,g12425);
  not NOT_4488(g13406,II20517);
  not NOT_4489(II20520,g13246);
  not NOT_4490(g13407,II20520);
  not NOT_4491(II20523,g13317);
  not NOT_4492(g13408,II20523);
  not NOT_4493(II20526,g12519);
  not NOT_4494(g13409,II20526);
  not NOT_4495(II20529,g13319);
  not NOT_4496(g13410,II20529);
  not NOT_4497(II20532,g13339);
  not NOT_4498(g13411,II20532);
  not NOT_4499(II20535,g13359);
  not NOT_4500(g13412,II20535);
  not NOT_4501(II20538,g13384);
  not NOT_4502(g13413,II20538);
  not NOT_4503(II20541,g11599);
  not NOT_4504(g13414,II20541);
  not NOT_4505(II20544,g11628);
  not NOT_4506(g13415,II20544);
  not NOT_4507(II20547,g13248);
  not NOT_4508(g13416,II20547);
  not NOT_4509(II20550,g13267);
  not NOT_4510(g13417,II20550);
  not NOT_4511(II20553,g13290);
  not NOT_4512(g13418,II20553);
  not NOT_4513(II20556,g12435);
  not NOT_4514(g13419,II20556);
  not NOT_4515(II20559,g11937);
  not NOT_4516(g13420,II20559);
  not NOT_4517(II20562,g11786);
  not NOT_4518(g13421,II20562);
  not NOT_4519(II20565,g12432);
  not NOT_4520(g13422,II20565);
  not NOT_4521(II20568,g13269);
  not NOT_4522(g13423,II20568);
  not NOT_4523(II20571,g13341);
  not NOT_4524(g13424,II20571);
  not NOT_4525(II20574,g12534);
  not NOT_4526(g13425,II20574);
  not NOT_4527(II20577,g13342);
  not NOT_4528(g13426,II20577);
  not NOT_4529(II20580,g13364);
  not NOT_4530(g13427,II20580);
  not NOT_4531(II20583,g13389);
  not NOT_4532(g13428,II20583);
  not NOT_4533(II20586,g11606);
  not NOT_4534(g13429,II20586);
  not NOT_4535(II20589,g11629);
  not NOT_4536(g13430,II20589);
  not NOT_4537(II20592,g11651);
  not NOT_4538(g13431,II20592);
  not NOT_4539(II20595,g13271);
  not NOT_4540(g13432,II20595);
  not NOT_4541(II20598,g13292);
  not NOT_4542(g13433,II20598);
  not NOT_4543(II20601,g13321);
  not NOT_4544(g13434,II20601);
  not NOT_4545(II20604,g12440);
  not NOT_4546(g13435,II20604);
  not NOT_4547(II20607,g11990);
  not NOT_4548(g13436,II20607);
  not NOT_4549(II20610,g11812);
  not NOT_4550(g13437,II20610);
  not NOT_4551(II20613,g12437);
  not NOT_4552(g13438,II20613);
  not NOT_4553(II20616,g13294);
  not NOT_4554(g13439,II20616);
  not NOT_4555(II20619,g13366);
  not NOT_4556(g13440,II20619);
  not NOT_4557(II20622,g12543);
  not NOT_4558(g13441,II20622);
  not NOT_4559(II20625,g13367);
  not NOT_4560(g13442,II20625);
  not NOT_4561(II20628,g13394);
  not NOT_4562(g13443,II20628);
  not NOT_4563(II20631,g11611);
  not NOT_4564(g13444,II20631);
  not NOT_4565(II20634,g11636);
  not NOT_4566(g13445,II20634);
  not NOT_4567(II20637,g11652);
  not NOT_4568(g13446,II20637);
  not NOT_4569(II20640,g11670);
  not NOT_4570(g13447,II20640);
  not NOT_4571(II20643,g13296);
  not NOT_4572(g13448,II20643);
  not NOT_4573(II20646,g13323);
  not NOT_4574(g13449,II20646);
  not NOT_4575(II20649,g13344);
  not NOT_4576(g13450,II20649);
  not NOT_4577(II20652,g12445);
  not NOT_4578(g13451,II20652);
  not NOT_4579(II20655,g12059);
  not NOT_4580(g13452,II20655);
  not NOT_4581(II20658,g11845);
  not NOT_4582(g13453,II20658);
  not NOT_4583(II20661,g12442);
  not NOT_4584(g13454,II20661);
  not NOT_4585(II20664,g13325);
  not NOT_4586(g13455,II20664);
  not NOT_4587(II20667,g13396);
  not NOT_4588(g13456,II20667);
  not NOT_4589(II20670,g12552);
  not NOT_4590(g13457,II20670);
  not NOT_4591(II20673,g13397);
  not NOT_4592(g13458,II20673);
  not NOT_4593(II20676,g11616);
  not NOT_4594(g13459,II20676);
  not NOT_4595(II20679,g11641);
  not NOT_4596(g13460,II20679);
  not NOT_4597(II20682,g11659);
  not NOT_4598(g13461,II20682);
  not NOT_4599(II20685,g11671);
  not NOT_4600(g13462,II20685);
  not NOT_4601(II20688,g11682);
  not NOT_4602(g13463,II20688);
  not NOT_4603(II20691,g13327);
  not NOT_4604(g13464,II20691);
  not NOT_4605(II20694,g13346);
  not NOT_4606(g13465,II20694);
  not NOT_4607(II20697,g13369);
  not NOT_4608(g13466,II20697);
  not NOT_4609(II20700,g12450);
  not NOT_4610(g13467,II20700);
  not NOT_4611(II20703,g12123);
  not NOT_4612(g13468,II20703);
  not NOT_4613(II20706,g11490);
  not NOT_4614(g13469,II20706);
  not NOT_4615(II20709,g13070);
  not NOT_4616(g13475,II20709);
  not NOT_4617(g13519,g13228);
  not NOT_4618(g13530,g13251);
  not NOT_4619(g13541,g13274);
  not NOT_4620(g13552,g13299);
  not NOT_4621(g13565,g12192);
  not NOT_4622(g13568,g11627);
  not NOT_4623(II20791,g13149);
  not NOT_4624(g13571,II20791);
  not NOT_4625(II20794,g13111);
  not NOT_4626(g13572,II20794);
  not NOT_4627(g13573,g12247);
  not NOT_4628(g13576,g11650);
  not NOT_4629(II20799,g13155);
  not NOT_4630(g13579,II20799);
  not NOT_4631(II20802,g13160);
  not NOT_4632(g13580,II20802);
  not NOT_4633(II20805,g13124);
  not NOT_4634(g13581,II20805);
  not NOT_4635(g13582,g12290);
  not NOT_4636(g13585,g11669);
  not NOT_4637(II20810,g13164);
  not NOT_4638(g13588,II20810);
  not NOT_4639(II20813,g13265);
  not NOT_4640(g13589,II20813);
  not NOT_4641(II20816,g12487);
  not NOT_4642(g13598,II20816);
  not NOT_4643(II20820,g13171);
  not NOT_4644(g13600,II20820);
  not NOT_4645(II20823,g13135);
  not NOT_4646(g13601,II20823);
  not NOT_4647(g13602,g12326);
  not NOT_4648(g13605,g11681);
  not NOT_4649(II20828,g13175);
  not NOT_4650(g13608,II20828);
  not NOT_4651(II20832,g12507);
  not NOT_4652(g13610,II20832);
  not NOT_4653(II20836,g13182);
  not NOT_4654(g13612,II20836);
  not NOT_4655(II20839,g13143);
  not NOT_4656(g13613,II20839);
  not NOT_4657(g13614,g11690);
  not NOT_4658(II20844,g12524);
  not NOT_4659(g13620,II20844);
  not NOT_4660(II20848,g13194);
  not NOT_4661(g13622,II20848);
  not NOT_4662(II20852,g12457);
  not NOT_4663(g13624,II20852);
  not NOT_4664(g13626,g11697);
  not NOT_4665(II20858,g12539);
  not NOT_4666(g13632,II20858);
  not NOT_4667(II20863,g12467);
  not NOT_4668(g13635,II20863);
  not NOT_4669(g13637,g11703);
  not NOT_4670(g13644,g13215);
  not NOT_4671(II20873,g12482);
  not NOT_4672(g13647,II20873);
  not NOT_4673(g13649,g11711);
  not NOT_4674(g13657,g12452);
  not NOT_4675(g13669,g13229);
  not NOT_4676(g13670,g13234);
  not NOT_4677(II20886,g12499);
  not NOT_4678(g13673,II20886);
  not NOT_4679(g13677,g12447);
  not NOT_4680(g13687,g12460);
  not NOT_4681(g13699,g13252);
  not NOT_4682(g13700,g13257);
  not NOT_4683(g13706,g12443);
  not NOT_4684(g13714,g12453);
  not NOT_4685(g13724,g12470);
  not NOT_4686(g13736,g13275);
  not NOT_4687(g13737,g13280);
  not NOT_4688(II20909,g13055);
  not NOT_4689(g13741,II20909);
  not NOT_4690(g13750,g12439);
  not NOT_4691(g13756,g12448);
  not NOT_4692(g13764,g12461);
  not NOT_4693(g13774,g12485);
  not NOT_4694(g13786,g13300);
  not NOT_4695(g13791,g12444);
  not NOT_4696(g13797,g12454);
  not NOT_4697(g13805,g12471);
  not NOT_4698(g13817,g13336);
  not NOT_4699(g13819,g12449);
  not NOT_4700(g13825,g12462);
  not NOT_4701(g13836,g13356);
  not NOT_4702(g13838,g13361);
  not NOT_4703(g13840,g12455);
  not NOT_4704(g13848,g11744);
  not NOT_4705(g13849,g13381);
  not NOT_4706(g13850,g13386);
  not NOT_4707(g13852,g13391);
  not NOT_4708(g13856,g11759);
  not NOT_4709(g13857,g11760);
  not NOT_4710(g13858,g11603);
  not NOT_4711(g13859,g11608);
  not NOT_4712(g13861,g11613);
  not NOT_4713(II20959,g11713);
  not NOT_4714(g13863,II20959);
  not NOT_4715(g13864,g11767);
  not NOT_4716(g13866,g11772);
  not NOT_4717(g13867,g11773);
  not NOT_4718(g13868,g11633);
  not NOT_4719(g13869,g11638);
  not NOT_4720(g13872,g11780);
  not NOT_4721(g13873,g12698);
  not NOT_4722(g13879,g11784);
  not NOT_4723(g13881,g11789);
  not NOT_4724(g13882,g11790);
  not NOT_4725(g13883,g11656);
  not NOT_4726(g13885,g11799);
  not NOT_4727(g13886,g12747);
  not NOT_4728(g13894,g11806);
  not NOT_4729(g13895,g12755);
  not NOT_4730(g13901,g11810);
  not NOT_4731(g13903,g11815);
  not NOT_4732(g13906,g11822);
  not NOT_4733(g13907,g12781);
  not NOT_4734(g13918,g11830);
  not NOT_4735(g13922,g11831);
  not NOT_4736(g13926,g11832);
  not NOT_4737(g13927,g12789);
  not NOT_4738(g13935,g11839);
  not NOT_4739(g13936,g12797);
  not NOT_4740(g13942,g11843);
  not NOT_4741(g13945,g11855);
  not NOT_4742(g13946,g12814);
  not NOT_4743(II21012,g12503);
  not NOT_4744(g13954,II21012);
  not NOT_4745(g13958,g11863);
  not NOT_4746(g13962,g11864);
  not NOT_4747(g13963,g12820);
  not NOT_4748(g13974,g11872);
  not NOT_4749(g13978,g11873);
  not NOT_4750(g13982,g11874);
  not NOT_4751(g13983,g12828);
  not NOT_4752(g13991,g11881);
  not NOT_4753(g13992,g12836);
  not NOT_4754(g13999,g11889);
  not NOT_4755(g14000,g11890);
  not NOT_4756(g14001,g12849);
  not NOT_4757(II21037,g12486);
  not NOT_4758(g14008,II21037);
  not NOT_4759(g14011,g11896);
  not NOT_4760(g14015,g11897);
  not NOT_4761(g14016,g12852);
  not NOT_4762(II21045,g12520);
  not NOT_4763(g14024,II21045);
  not NOT_4764(g14028,g11905);
  not NOT_4765(g14032,g11906);
  not NOT_4766(g14033,g12858);
  not NOT_4767(g14044,g11914);
  not NOT_4768(g14048,g11915);
  not NOT_4769(g14052,g11916);
  not NOT_4770(g14053,g12866);
  not NOT_4771(g14061,g11928);
  not NOT_4772(g14062,g12880);
  not NOT_4773(II21064,g13147);
  not NOT_4774(g14068,II21064);
  not NOT_4775(g14071,g11934);
  not NOT_4776(g14079,g11935);
  not NOT_4777(g14086,g11938);
  not NOT_4778(g14090,g11939);
  not NOT_4779(g14091,g11940);
  not NOT_4780(g14092,g12890);
  not NOT_4781(II21075,g12506);
  not NOT_4782(g14099,II21075);
  not NOT_4783(g14102,g11946);
  not NOT_4784(g14106,g11947);
  not NOT_4785(g14107,g12893);
  not NOT_4786(II21083,g12535);
  not NOT_4787(g14115,II21083);
  not NOT_4788(g14119,g11955);
  not NOT_4789(g14123,g11956);
  not NOT_4790(g14124,g12899);
  not NOT_4791(g14135,g11964);
  not NOT_4792(g14139,g11965);
  not NOT_4793(II21096,g11749);
  not NOT_4794(g14144,II21096);
  not NOT_4795(g14148,g12912);
  not NOT_4796(g14153,g12913);
  not NOT_4797(g14158,g11974);
  not NOT_4798(g14165,g11975);
  not NOT_4799(g14171,g11979);
  not NOT_4800(g14175,g11980);
  not NOT_4801(g14176,g11981);
  not NOT_4802(g14177,g12920);
  not NOT_4803(II21108,g13150);
  not NOT_4804(g14183,II21108);
  not NOT_4805(g14186,g11987);
  not NOT_4806(g14194,g11988);
  not NOT_4807(g14201,g11991);
  not NOT_4808(g14205,g11992);
  not NOT_4809(g14206,g11993);
  not NOT_4810(g14207,g12930);
  not NOT_4811(II21119,g12523);
  not NOT_4812(g14214,II21119);
  not NOT_4813(g14217,g11999);
  not NOT_4814(g14221,g12000);
  not NOT_4815(g14222,g12933);
  not NOT_4816(II21127,g12544);
  not NOT_4817(g14230,II21127);
  not NOT_4818(g14234,g12008);
  not NOT_4819(g14238,g12939);
  not NOT_4820(g14244,g12026);
  not NOT_4821(g14249,g12034);
  not NOT_4822(g14252,g12035);
  not NOT_4823(g14256,g12036);
  not NOT_4824(II21137,g11749);
  not NOT_4825(g14259,II21137);
  not NOT_4826(g14263,g12941);
  not NOT_4827(g14268,g12942);
  not NOT_4828(g14273,g12043);
  not NOT_4829(g14280,g12044);
  not NOT_4830(g14286,g12048);
  not NOT_4831(g14290,g12049);
  not NOT_4832(g14291,g12050);
  not NOT_4833(g14292,g12949);
  not NOT_4834(II21149,g13156);
  not NOT_4835(g14298,II21149);
  not NOT_4836(g14301,g12056);
  not NOT_4837(g14309,g12057);
  not NOT_4838(g14316,g12060);
  not NOT_4839(g14320,g12061);
  not NOT_4840(g14321,g12062);
  not NOT_4841(g14322,g12959);
  not NOT_4842(II21160,g12538);
  not NOT_4843(g14329,II21160);
  not NOT_4844(g14332,g12068);
  not NOT_4845(II21165,g13110);
  not NOT_4846(g14337,II21165);
  not NOT_4847(g14342,g12967);
  not NOT_4848(g14347,g12079);
  not NOT_4849(g14352,g12081);
  not NOT_4850(g14355,g12082);
  not NOT_4851(g14359,g12083);
  not NOT_4852(g14360,g12968);
  not NOT_4853(g14366,g12090);
  not NOT_4854(g14371,g12098);
  not NOT_4855(g14374,g12099);
  not NOT_4856(g14378,g12100);
  not NOT_4857(II21178,g11749);
  not NOT_4858(g14381,II21178);
  not NOT_4859(g14385,g12970);
  not NOT_4860(g14390,g12971);
  not NOT_4861(g14395,g12107);
  not NOT_4862(g14402,g12108);
  not NOT_4863(g14408,g12112);
  not NOT_4864(g14412,g12113);
  not NOT_4865(g14413,g12114);
  not NOT_4866(g14414,g12978);
  not NOT_4867(II21190,g13165);
  not NOT_4868(g14420,II21190);
  not NOT_4869(g14423,g12120);
  not NOT_4870(g14431,g12121);
  not NOT_4871(g14438,g12124);
  not NOT_4872(g14442,g11768);
  not NOT_4873(g14450,g12146);
  not NOT_4874(g14454,g12991);
  not NOT_4875(g14459,g12151);
  not NOT_4876(g14464,g12153);
  not NOT_4877(g14467,g12154);
  not NOT_4878(g14471,g12155);
  not NOT_4879(g14472,g12992);
  not NOT_4880(g14478,g12162);
  not NOT_4881(g14483,g12170);
  not NOT_4882(g14486,g12171);
  not NOT_4883(g14490,g12172);
  not NOT_4884(II21208,g11749);
  not NOT_4885(g14493,II21208);
  not NOT_4886(g14497,g12994);
  not NOT_4887(g14502,g12995);
  not NOT_4888(g14507,g12179);
  not NOT_4889(g14514,g12180);
  not NOT_4890(g14520,g12184);
  not NOT_4891(g14524,g12185);
  not NOT_4892(g14525,g12195);
  not NOT_4893(g14529,g11785);
  not NOT_4894(g14537,g12208);
  not NOT_4895(g14541,g13001);
  not NOT_4896(g14546,g12213);
  not NOT_4897(g14551,g12215);
  not NOT_4898(g14554,g12216);
  not NOT_4899(g14558,g12217);
  not NOT_4900(g14559,g13002);
  not NOT_4901(g14565,g12224);
  not NOT_4902(g14570,g12232);
  not NOT_4903(g14573,g12233);
  not NOT_4904(g14577,g12234);
  not NOT_4905(g14580,g12250);
  not NOT_4906(g14584,g11811);
  not NOT_4907(g14592,g12263);
  not NOT_4908(g14596,g13022);
  not NOT_4909(g14601,g12268);
  not NOT_4910(g14606,g12270);
  not NOT_4911(g14609,g12271);
  not NOT_4912(g14613,g12272);
  not NOT_4913(g14614,g12293);
  not NOT_4914(g14618,g11844);
  not NOT_4915(g14626,g12306);
  not NOT_4916(II21241,g13378);
  not NOT_4917(g14630,II21241);
  not NOT_4918(g14637,g12329);
  not NOT_4919(g14641,g11823);
  not NOT_4920(II21246,g11624);
  not NOT_4921(g14642,II21246);
  not NOT_4922(II21249,g11600);
  not NOT_4923(g14650,II21249);
  not NOT_4924(II21252,g11644);
  not NOT_4925(g14657,II21252);
  not NOT_4926(g14668,g11865);
  not NOT_4927(II21256,g11647);
  not NOT_4928(g14669,II21256);
  not NOT_4929(II21259,g11630);
  not NOT_4930(g14677,II21259);
  not NOT_4931(II21262,g11713);
  not NOT_4932(g14684,II21262);
  not NOT_4933(g14685,g12245);
  not NOT_4934(II21267,g11663);
  not NOT_4935(g14691,II21267);
  not NOT_4936(g14702,g11907);
  not NOT_4937(II21271,g11666);
  not NOT_4938(g14703,II21271);
  not NOT_4939(II21274,g11653);
  not NOT_4940(g14711,II21274);
  not NOT_4941(II21277,g12430);
  not NOT_4942(g14718,II21277);
  not NOT_4943(g14719,g12288);
  not NOT_4944(II21282,g11675);
  not NOT_4945(g14725,II21282);
  not NOT_4946(g14736,g11957);
  not NOT_4947(II21286,g11678);
  not NOT_4948(g14737,II21286);
  not NOT_4949(II21289,g12434);
  not NOT_4950(g14745,II21289);
  not NOT_4951(II21292,g11888);
  not NOT_4952(g14746,II21292);
  not NOT_4953(g14747,g12324);
  not NOT_4954(II21297,g11687);
  not NOT_4955(g14753,II21297);
  not NOT_4956(g14764,g11791);
  not NOT_4957(II21301,g12438);
  not NOT_4958(g14765,II21301);
  not NOT_4959(II21304,g11927);
  not NOT_4960(g14766,II21304);
  not NOT_4961(g14768,g12352);
  not NOT_4962(II21310,g12332);
  not NOT_4963(g14774,II21310);
  not NOT_4964(II21313,g11743);
  not NOT_4965(g14775,II21313);
  not NOT_4966(g14776,g12033);
  not NOT_4967(g14794,g11848);
  not NOT_4968(II21318,g12362);
  not NOT_4969(g14795,II21318);
  not NOT_4970(II21321,g11758);
  not NOT_4971(g14796,II21321);
  not NOT_4972(g14797,g12080);
  not NOT_4973(g14811,g12097);
  not NOT_4974(II21326,g12378);
  not NOT_4975(g14829,II21326);
  not NOT_4976(II21329,g11766);
  not NOT_4977(g14830,II21329);
  not NOT_4978(g14831,g11828);
  not NOT_4979(g14837,g12145);
  not NOT_4980(g14849,g12152);
  not NOT_4981(g14863,g12169);
  not NOT_4982(g14881,g11923);
  not NOT_4983(II21337,g12408);
  not NOT_4984(g14882,II21337);
  not NOT_4985(II21340,g11779);
  not NOT_4986(g14883,II21340);
  not NOT_4987(g14885,g11860);
  not NOT_4988(g14895,g12193);
  not NOT_4989(g14904,g11870);
  not NOT_4990(g14910,g12207);
  not NOT_4991(g14922,g12214);
  not NOT_4992(g14936,g12231);
  not NOT_4993(II21351,g12420);
  not NOT_4994(g14954,II21351);
  not NOT_4995(II21354,g11798);
  not NOT_4996(g14955,II21354);
  not NOT_4997(g14959,g11976);
  not NOT_4998(II21361,g13026);
  not NOT_4999(g14960,II21361);
  not NOT_5000(II21364,g13028);
  not NOT_5001(g14963,II21364);
  not NOT_5002(g14966,g11902);
  not NOT_5003(g14976,g12248);
  not NOT_5004(g14985,g11912);
  not NOT_5005(g14991,g12262);
  not NOT_5006(g15003,g12269);
  not NOT_5007(g15017,g12009);
  not NOT_5008(II21374,g12424);
  not NOT_5009(g15018,II21374);
  not NOT_5010(II21377,g11821);
  not NOT_5011(g15019,II21377);
  not NOT_5012(II21381,g13157);
  not NOT_5013(g15021,II21381);
  not NOT_5014(g15022,g11781);
  not NOT_5015(g15032,g12027);
  not NOT_5016(g15033,g12030);
  not NOT_5017(II21389,g12883);
  not NOT_5018(g15034,II21389);
  not NOT_5019(II21392,g13020);
  not NOT_5020(g15037,II21392);
  not NOT_5021(II21395,g13034);
  not NOT_5022(g15040,II21395);
  not NOT_5023(II21398,g13021);
  not NOT_5024(g15043,II21398);
  not NOT_5025(g15048,g12045);
  not NOT_5026(II21404,g13037);
  not NOT_5027(g15049,II21404);
  not NOT_5028(II21407,g13039);
  not NOT_5029(g15052,II21407);
  not NOT_5030(g15055,g11952);
  not NOT_5031(g15065,g12291);
  not NOT_5032(g15074,g11962);
  not NOT_5033(g15080,g12305);
  not NOT_5034(II21415,g11854);
  not NOT_5035(g15092,II21415);
  not NOT_5036(II21420,g13166);
  not NOT_5037(g15095,II21420);
  not NOT_5038(g15096,g11800);
  not NOT_5039(II21426,g11661);
  not NOT_5040(g15106,II21426);
  not NOT_5041(II21429,g13027);
  not NOT_5042(g15109,II21429);
  not NOT_5043(II21432,g13044);
  not NOT_5044(g15112,II21432);
  not NOT_5045(II21435,g11662);
  not NOT_5046(g15115,II21435);
  not NOT_5047(g15118,g11807);
  not NOT_5048(g15128,g12091);
  not NOT_5049(g15129,g12094);
  not NOT_5050(II21443,g12923);
  not NOT_5051(g15130,II21443);
  not NOT_5052(II21446,g13029);
  not NOT_5053(g15133,II21446);
  not NOT_5054(II21449,g13047);
  not NOT_5055(g15136,II21449);
  not NOT_5056(II21452,g13030);
  not NOT_5057(g15139,II21452);
  not NOT_5058(g15144,g12109);
  not NOT_5059(II21458,g13050);
  not NOT_5060(g15145,II21458);
  not NOT_5061(II21461,g13052);
  not NOT_5062(g15148,II21461);
  not NOT_5063(g15151,g12005);
  not NOT_5064(g15161,g12327);
  not NOT_5065(g15170,g12125);
  not NOT_5066(g15174,g12136);
  not NOT_5067(g15175,g12139);
  not NOT_5068(g15176,g12142);
  not NOT_5069(g15177,g12339);
  not NOT_5070(II21476,g11672);
  not NOT_5071(g15179,II21476);
  not NOT_5072(II21479,g13035);
  not NOT_5073(g15182,II21479);
  not NOT_5074(II21482,g13058);
  not NOT_5075(g15185,II21482);
  not NOT_5076(g15188,g11833);
  not NOT_5077(II21488,g11673);
  not NOT_5078(g15198,II21488);
  not NOT_5079(II21491,g13038);
  not NOT_5080(g15201,II21491);
  not NOT_5081(II21494,g13061);
  not NOT_5082(g15204,II21494);
  not NOT_5083(II21497,g11674);
  not NOT_5084(g15207,II21497);
  not NOT_5085(g15210,g11840);
  not NOT_5086(g15220,g12163);
  not NOT_5087(g15221,g12166);
  not NOT_5088(II21505,g12952);
  not NOT_5089(g15222,II21505);
  not NOT_5090(II21508,g13040);
  not NOT_5091(g15225,II21508);
  not NOT_5092(II21511,g13064);
  not NOT_5093(g15228,II21511);
  not NOT_5094(II21514,g13041);
  not NOT_5095(g15231,II21514);
  not NOT_5096(g15236,g12181);
  not NOT_5097(II21520,g13067);
  not NOT_5098(g15237,II21520);
  not NOT_5099(II21523,g13069);
  not NOT_5100(g15240,II21523);
  not NOT_5101(II21531,g11683);
  not NOT_5102(g15248,II21531);
  not NOT_5103(II21534,g13045);
  not NOT_5104(g15251,II21534);
  not NOT_5105(II21537,g13071);
  not NOT_5106(g15254,II21537);
  not NOT_5107(g15260,g12198);
  not NOT_5108(g15261,g12201);
  not NOT_5109(g15262,g12204);
  not NOT_5110(g15263,g12369);
  not NOT_5111(II21548,g11684);
  not NOT_5112(g15265,II21548);
  not NOT_5113(II21551,g13048);
  not NOT_5114(g15268,II21551);
  not NOT_5115(II21554,g13074);
  not NOT_5116(g15271,II21554);
  not NOT_5117(g15274,g11875);
  not NOT_5118(II21560,g11685);
  not NOT_5119(g15284,II21560);
  not NOT_5120(II21563,g13051);
  not NOT_5121(g15287,II21563);
  not NOT_5122(II21566,g13077);
  not NOT_5123(g15290,II21566);
  not NOT_5124(II21569,g11686);
  not NOT_5125(g15293,II21569);
  not NOT_5126(g15296,g11882);
  not NOT_5127(g15306,g12225);
  not NOT_5128(g15307,g12228);
  not NOT_5129(II21577,g12981);
  not NOT_5130(g15308,II21577);
  not NOT_5131(II21580,g13053);
  not NOT_5132(g15311,II21580);
  not NOT_5133(II21583,g13080);
  not NOT_5134(g15314,II21583);
  not NOT_5135(II21586,g13054);
  not NOT_5136(g15317,II21586);
  not NOT_5137(g15322,g12239);
  not NOT_5138(g15323,g12242);
  not NOT_5139(II21595,g11691);
  not NOT_5140(g15326,II21595);
  not NOT_5141(II21598,g13059);
  not NOT_5142(g15329,II21598);
  not NOT_5143(II21601,g13087);
  not NOT_5144(g15332,II21601);
  not NOT_5145(II21609,g11692);
  not NOT_5146(g15340,II21609);
  not NOT_5147(II21612,g13062);
  not NOT_5148(g15343,II21612);
  not NOT_5149(II21615,g13090);
  not NOT_5150(g15346,II21615);
  not NOT_5151(g15352,g12253);
  not NOT_5152(g15353,g12256);
  not NOT_5153(g15354,g12259);
  not NOT_5154(g15355,g12388);
  not NOT_5155(II21626,g11693);
  not NOT_5156(g15357,II21626);
  not NOT_5157(II21629,g13065);
  not NOT_5158(g15360,II21629);
  not NOT_5159(II21632,g13093);
  not NOT_5160(g15363,II21632);
  not NOT_5161(g15366,g11917);
  not NOT_5162(II21638,g11694);
  not NOT_5163(g15376,II21638);
  not NOT_5164(II21641,g13068);
  not NOT_5165(g15379,II21641);
  not NOT_5166(II21644,g13096);
  not NOT_5167(g15382,II21644);
  not NOT_5168(II21647,g11695);
  not NOT_5169(g15385,II21647);
  not NOT_5170(g15390,g12279);
  not NOT_5171(II21655,g11696);
  not NOT_5172(g15393,II21655);
  not NOT_5173(II21658,g13072);
  not NOT_5174(g15396,II21658);
  not NOT_5175(II21661,g13098);
  not NOT_5176(g15399,II21661);
  not NOT_5177(II21666,g13100);
  not NOT_5178(g15404,II21666);
  not NOT_5179(g15408,g12282);
  not NOT_5180(g15409,g12285);
  not NOT_5181(II21674,g11698);
  not NOT_5182(g15412,II21674);
  not NOT_5183(II21677,g13075);
  not NOT_5184(g15415,II21677);
  not NOT_5185(II21680,g13102);
  not NOT_5186(g15418,II21680);
  not NOT_5187(II21688,g11699);
  not NOT_5188(g15426,II21688);
  not NOT_5189(II21691,g13078);
  not NOT_5190(g15429,II21691);
  not NOT_5191(II21694,g13105);
  not NOT_5192(g15432,II21694);
  not NOT_5193(g15438,g12296);
  not NOT_5194(g15439,g12299);
  not NOT_5195(g15440,g12302);
  not NOT_5196(g15441,g12418);
  not NOT_5197(II21705,g11700);
  not NOT_5198(g15443,II21705);
  not NOT_5199(II21708,g13081);
  not NOT_5200(g15446,II21708);
  not NOT_5201(II21711,g13108);
  not NOT_5202(g15449,II21711);
  not NOT_5203(g15458,g12312);
  not NOT_5204(II21720,g11701);
  not NOT_5205(g15461,II21720);
  not NOT_5206(II21723,g13088);
  not NOT_5207(g15464,II21723);
  not NOT_5208(II21726,g13112);
  not NOT_5209(g15467,II21726);
  not NOT_5210(II21730,g13089);
  not NOT_5211(g15471,II21730);
  not NOT_5212(g15474,g12315);
  not NOT_5213(II21736,g11702);
  not NOT_5214(g15477,II21736);
  not NOT_5215(II21739,g13091);
  not NOT_5216(g15480,II21739);
  not NOT_5217(II21742,g13114);
  not NOT_5218(g15483,II21742);
  not NOT_5219(II21747,g13116);
  not NOT_5220(g15488,II21747);
  not NOT_5221(g15492,g12318);
  not NOT_5222(g15493,g12321);
  not NOT_5223(II21755,g11704);
  not NOT_5224(g15496,II21755);
  not NOT_5225(II21758,g13094);
  not NOT_5226(g15499,II21758);
  not NOT_5227(II21761,g13118);
  not NOT_5228(g15502,II21761);
  not NOT_5229(II21769,g11705);
  not NOT_5230(g15510,II21769);
  not NOT_5231(II21772,g13097);
  not NOT_5232(g15513,II21772);
  not NOT_5233(II21775,g13121);
  not NOT_5234(g15516,II21775);
  not NOT_5235(II21780,g13305);
  not NOT_5236(g15521,II21780);
  not NOT_5237(g15524,g12333);
  not NOT_5238(g15525,g12336);
  not NOT_5239(II21787,g11707);
  not NOT_5240(g15528,II21787);
  not NOT_5241(II21790,g13099);
  not NOT_5242(g15531,II21790);
  not NOT_5243(II21793,g13123);
  not NOT_5244(g15534,II21793);
  not NOT_5245(II21796,g11708);
  not NOT_5246(g15537,II21796);
  not NOT_5247(g15544,g12340);
  not NOT_5248(II21803,g11709);
  not NOT_5249(g15547,II21803);
  not NOT_5250(II21806,g13103);
  not NOT_5251(g15550,II21806);
  not NOT_5252(II21809,g13125);
  not NOT_5253(g15553,II21809);
  not NOT_5254(II21813,g13104);
  not NOT_5255(g15557,II21813);
  not NOT_5256(g15560,g12343);
  not NOT_5257(II21819,g11710);
  not NOT_5258(g15563,II21819);
  not NOT_5259(II21822,g13106);
  not NOT_5260(g15566,II21822);
  not NOT_5261(II21825,g13127);
  not NOT_5262(g15569,II21825);
  not NOT_5263(II21830,g13129);
  not NOT_5264(g15574,II21830);
  not NOT_5265(g15578,g12346);
  not NOT_5266(g15579,g12349);
  not NOT_5267(II21838,g11712);
  not NOT_5268(g15582,II21838);
  not NOT_5269(II21841,g13109);
  not NOT_5270(g15585,II21841);
  not NOT_5271(II21844,g13131);
  not NOT_5272(g15588,II21844);
  not NOT_5273(II21852,g11716);
  not NOT_5274(g15596,II21852);
  not NOT_5275(II21855,g13113);
  not NOT_5276(g15599,II21855);
  not NOT_5277(g15602,g12363);
  not NOT_5278(g15603,g12366);
  not NOT_5279(II21862,g11717);
  not NOT_5280(g15606,II21862);
  not NOT_5281(II21865,g13115);
  not NOT_5282(g15609,II21865);
  not NOT_5283(II21868,g13134);
  not NOT_5284(g15612,II21868);
  not NOT_5285(II21871,g11718);
  not NOT_5286(g15615,II21871);
  not NOT_5287(g15622,g12370);
  not NOT_5288(II21878,g11719);
  not NOT_5289(g15625,II21878);
  not NOT_5290(II21881,g13119);
  not NOT_5291(g15628,II21881);
  not NOT_5292(II21884,g13136);
  not NOT_5293(g15631,II21884);
  not NOT_5294(II21888,g13120);
  not NOT_5295(g15635,II21888);
  not NOT_5296(g15638,g12373);
  not NOT_5297(II21894,g11720);
  not NOT_5298(g15641,II21894);
  not NOT_5299(II21897,g13122);
  not NOT_5300(g15644,II21897);
  not NOT_5301(II21900,g13138);
  not NOT_5302(g15647,II21900);
  not NOT_5303(II21905,g13140);
  not NOT_5304(g15652,II21905);
  not NOT_5305(II21908,g13082);
  not NOT_5306(g15655,II21908);
  not NOT_5307(g15659,g11706);
  not NOT_5308(g15665,g12379);
  not NOT_5309(II21918,g11721);
  not NOT_5310(g15667,II21918);
  not NOT_5311(II21923,g11722);
  not NOT_5312(g15672,II21923);
  not NOT_5313(II21926,g13126);
  not NOT_5314(g15675,II21926);
  not NOT_5315(g15678,g12382);
  not NOT_5316(g15679,g12385);
  not NOT_5317(II21933,g11723);
  not NOT_5318(g15682,II21933);
  not NOT_5319(II21936,g13128);
  not NOT_5320(g15685,II21936);
  not NOT_5321(II21939,g13142);
  not NOT_5322(g15688,II21939);
  not NOT_5323(II21942,g11724);
  not NOT_5324(g15691,II21942);
  not NOT_5325(g15698,g12389);
  not NOT_5326(II21949,g11725);
  not NOT_5327(g15701,II21949);
  not NOT_5328(II21952,g13132);
  not NOT_5329(g15704,II21952);
  not NOT_5330(II21955,g13144);
  not NOT_5331(g15707,II21955);
  not NOT_5332(II21959,g13133);
  not NOT_5333(g15711,II21959);
  not NOT_5334(II21962,g13004);
  not NOT_5335(g15714,II21962);
  not NOT_5336(g15722,g13011);
  not NOT_5337(g15724,g12409);
  not NOT_5338(II21974,g11726);
  not NOT_5339(g15726,II21974);
  not NOT_5340(II21979,g11727);
  not NOT_5341(g15731,II21979);
  not NOT_5342(II21982,g13137);
  not NOT_5343(g15734,II21982);
  not NOT_5344(g15737,g12412);
  not NOT_5345(g15738,g12415);
  not NOT_5346(II21989,g11728);
  not NOT_5347(g15741,II21989);
  not NOT_5348(II21992,g13139);
  not NOT_5349(g15744,II21992);
  not NOT_5350(II21995,g13146);
  not NOT_5351(g15747,II21995);
  not NOT_5352(II21998,g11729);
  not NOT_5353(g15750,II21998);
  not NOT_5354(g15762,g13011);
  not NOT_5355(g15764,g12421);
  not NOT_5356(II22014,g11730);
  not NOT_5357(g15766,II22014);
  not NOT_5358(II22019,g11731);
  not NOT_5359(g15771,II22019);
  not NOT_5360(II22022,g13145);
  not NOT_5361(g15774,II22022);
  not NOT_5362(II22025,g11617);
  not NOT_5363(g15777,II22025);
  not NOT_5364(g15790,g13011);
  not NOT_5365(g15792,g12426);
  not NOT_5366(II22044,g11733);
  not NOT_5367(g15794,II22044);
  not NOT_5368(g15800,g12909);
  not NOT_5369(g15813,g13011);
  not NOT_5370(g15859,g13378);
  not NOT_5371(II22120,g12909);
  not NOT_5372(g15876,II22120);
  not NOT_5373(g15880,g11624);
  not NOT_5374(g15890,g11600);
  not NOT_5375(g15904,g11644);
  not NOT_5376(g15913,g11647);
  not NOT_5377(g15923,g11630);
  not NOT_5378(g15933,g11663);
  not NOT_5379(g15942,g11666);
  not NOT_5380(g15952,g11653);
  not NOT_5381(g15962,g11675);
  not NOT_5382(g15971,g11678);
  not NOT_5383(g15981,g11687);
  not NOT_5384(II22163,g12433);
  not NOT_5385(g15989,II22163);
  not NOT_5386(g15991,g12548);
  not NOT_5387(g15994,g12555);
  not NOT_5388(g15997,g12561);
  not NOT_5389(g16001,g12601);
  not NOT_5390(g16002,g12604);
  not NOT_5391(g16005,g12608);
  not NOT_5392(g16007,g12647);
  not NOT_5393(g16011,g12651);
  not NOT_5394(g16012,g12654);
  not NOT_5395(g16013,g12692);
  not NOT_5396(g16014,g12695);
  not NOT_5397(g16023,g12699);
  not NOT_5398(g16024,g12702);
  not NOT_5399(g16025,g12705);
  not NOT_5400(g16026,g12708);
  not NOT_5401(g16027,g12744);
  not NOT_5402(g16034,g12749);
  not NOT_5403(g16035,g12752);
  not NOT_5404(g16039,g12756);
  not NOT_5405(g16040,g12759);
  not NOT_5406(g16041,g12762);
  not NOT_5407(g16042,g12765);
  not NOT_5408(g16043,g12769);
  not NOT_5409(g16044,g12772);
  not NOT_5410(g16054,g12783);
  not NOT_5411(g16055,g12786);
  not NOT_5412(g16056,g12791);
  not NOT_5413(g16057,g12794);
  not NOT_5414(g16061,g12798);
  not NOT_5415(g16062,g12801);
  not NOT_5416(g16063,g12804);
  not NOT_5417(g16064,g12808);
  not NOT_5418(g16065,g12811);
  not NOT_5419(g16075,g11861);
  not NOT_5420(g16088,g12816);
  not NOT_5421(g16090,g12822);
  not NOT_5422(g16091,g12825);
  not NOT_5423(g16092,g12830);
  not NOT_5424(g16093,g12833);
  not NOT_5425(g16097,g12837);
  not NOT_5426(g16098,g12840);
  not NOT_5427(g16099,g12844);
  not NOT_5428(g16113,g11903);
  not NOT_5429(g16126,g12854);
  not NOT_5430(g16128,g12860);
  not NOT_5431(g16129,g12863);
  not NOT_5432(g16130,g12868);
  not NOT_5433(g16131,g12871);
  not NOT_5434(g16142,g13057);
  not NOT_5435(g16154,g12194);
  not NOT_5436(g16164,g11953);
  not NOT_5437(g16177,g12895);
  not NOT_5438(g16179,g12901);
  not NOT_5439(g16180,g12904);
  not NOT_5440(g16189,g13043);
  not NOT_5441(g16201,g13073);
  not NOT_5442(g16213,g12249);
  not NOT_5443(g16223,g12006);
  not NOT_5444(g16236,g12935);
  not NOT_5445(g16243,g13033);
  not NOT_5446(g16254,g13060);
  not NOT_5447(g16266,g13092);
  not NOT_5448(g16278,g12292);
  not NOT_5449(g16287,g12962);
  not NOT_5450(g16293,g13025);
  not NOT_5451(II22382,g520);
  not NOT_5452(g16297,II22382);
  not NOT_5453(g16302,g13046);
  not NOT_5454(g16313,g13076);
  not NOT_5455(g16325,g13107);
  not NOT_5456(g16337,g12328);
  not NOT_5457(g16351,g13036);
  not NOT_5458(II22414,g1206);
  not NOT_5459(g16355,II22414);
  not NOT_5460(g16360,g13063);
  not NOT_5461(g16371,g13095);
  not NOT_5462(g16395,g13049);
  not NOT_5463(II22444,g1900);
  not NOT_5464(g16399,II22444);
  not NOT_5465(g16404,g13079);
  not NOT_5466(g16433,g13066);
  not NOT_5467(II22475,g2594);
  not NOT_5468(g16437,II22475);
  not NOT_5469(g16466,g12017);
  not NOT_5470(II22503,g13598);
  not NOT_5471(g16467,II22503);
  not NOT_5472(II22506,g13624);
  not NOT_5473(g16468,II22506);
  not NOT_5474(II22509,g13610);
  not NOT_5475(g16469,II22509);
  not NOT_5476(II22512,g13635);
  not NOT_5477(g16470,II22512);
  not NOT_5478(II22515,g13620);
  not NOT_5479(g16471,II22515);
  not NOT_5480(II22518,g13647);
  not NOT_5481(g16472,II22518);
  not NOT_5482(II22521,g13632);
  not NOT_5483(g16473,II22521);
  not NOT_5484(II22524,g13673);
  not NOT_5485(g16474,II22524);
  not NOT_5486(II22527,g13469);
  not NOT_5487(g16475,II22527);
  not NOT_5488(II22530,g14774);
  not NOT_5489(g16476,II22530);
  not NOT_5490(II22533,g14795);
  not NOT_5491(g16477,II22533);
  not NOT_5492(II22536,g14829);
  not NOT_5493(g16478,II22536);
  not NOT_5494(II22539,g14882);
  not NOT_5495(g16479,II22539);
  not NOT_5496(II22542,g14954);
  not NOT_5497(g16480,II22542);
  not NOT_5498(II22545,g15018);
  not NOT_5499(g16481,II22545);
  not NOT_5500(II22548,g14718);
  not NOT_5501(g16482,II22548);
  not NOT_5502(II22551,g14745);
  not NOT_5503(g16483,II22551);
  not NOT_5504(II22554,g14765);
  not NOT_5505(g16484,II22554);
  not NOT_5506(II22557,g14775);
  not NOT_5507(g16485,II22557);
  not NOT_5508(II22560,g14796);
  not NOT_5509(g16486,II22560);
  not NOT_5510(II22563,g14830);
  not NOT_5511(g16487,II22563);
  not NOT_5512(II22566,g14883);
  not NOT_5513(g16488,II22566);
  not NOT_5514(II22569,g14955);
  not NOT_5515(g16489,II22569);
  not NOT_5516(II22572,g15019);
  not NOT_5517(g16490,II22572);
  not NOT_5518(II22575,g15092);
  not NOT_5519(g16491,II22575);
  not NOT_5520(II22578,g14746);
  not NOT_5521(g16492,II22578);
  not NOT_5522(II22581,g14766);
  not NOT_5523(g16493,II22581);
  not NOT_5524(II22584,g15989);
  not NOT_5525(g16494,II22584);
  not NOT_5526(II22587,g14684);
  not NOT_5527(g16495,II22587);
  not NOT_5528(II22590,g13863);
  not NOT_5529(g16496,II22590);
  not NOT_5530(II22593,g15876);
  not NOT_5531(g16497,II22593);
  not NOT_5532(g16501,g14158);
  not NOT_5533(II22599,g14966);
  not NOT_5534(g16506,II22599);
  not NOT_5535(g16507,g14186);
  not NOT_5536(II22604,g15080);
  not NOT_5537(g16514,II22604);
  not NOT_5538(g16515,g14244);
  not NOT_5539(g16523,g14273);
  not NOT_5540(II22611,g15055);
  not NOT_5541(g16528,II22611);
  not NOT_5542(g16529,g14301);
  not NOT_5543(II22618,g14630);
  not NOT_5544(g16540,II22618);
  not NOT_5545(g16543,g14347);
  not NOT_5546(g16546,g14366);
  not NOT_5547(g16554,g14395);
  not NOT_5548(II22626,g15151);
  not NOT_5549(g16559,II22626);
  not NOT_5550(g16560,g14423);
  not NOT_5551(II22640,g14650);
  not NOT_5552(g16572,II22640);
  not NOT_5553(g16575,g14459);
  not NOT_5554(g16578,g14478);
  not NOT_5555(g16586,g14507);
  not NOT_5556(II22651,g14677);
  not NOT_5557(g16596,II22651);
  not NOT_5558(g16599,g14546);
  not NOT_5559(g16602,g14565);
  not NOT_5560(II22657,g14657);
  not NOT_5561(g16608,II22657);
  not NOT_5562(II22663,g14711);
  not NOT_5563(g16616,II22663);
  not NOT_5564(g16619,g14601);
  not NOT_5565(II22667,g14642);
  not NOT_5566(g16622,II22667);
  not NOT_5567(II22671,g14691);
  not NOT_5568(g16626,II22671);
  not NOT_5569(II22676,g14630);
  not NOT_5570(g16633,II22676);
  not NOT_5571(II22679,g14669);
  not NOT_5572(g16636,II22679);
  not NOT_5573(II22683,g14725);
  not NOT_5574(g16640,II22683);
  not NOT_5575(II22687,g14650);
  not NOT_5576(g16644,II22687);
  not NOT_5577(II22690,g14703);
  not NOT_5578(g16647,II22690);
  not NOT_5579(II22694,g14753);
  not NOT_5580(g16651,II22694);
  not NOT_5581(II22699,g14677);
  not NOT_5582(g16656,II22699);
  not NOT_5583(II22702,g14737);
  not NOT_5584(g16659,II22702);
  not NOT_5585(g16665,g14776);
  not NOT_5586(II22715,g14711);
  not NOT_5587(g16673,II22715);
  not NOT_5588(II22718,g14657);
  not NOT_5589(g16676,II22718);
  not NOT_5590(g16682,g14797);
  not NOT_5591(g16686,g14811);
  not NOT_5592(II22726,g14642);
  not NOT_5593(g16694,II22726);
  not NOT_5594(g16697,g14837);
  not NOT_5595(II22730,g14691);
  not NOT_5596(g16702,II22730);
  not NOT_5597(g16708,g14849);
  not NOT_5598(g16712,g14863);
  not NOT_5599(II22737,g14630);
  not NOT_5600(g16719,II22737);
  not NOT_5601(g16722,g14895);
  not NOT_5602(II22741,g14669);
  not NOT_5603(g16725,II22741);
  not NOT_5604(g16728,g14910);
  not NOT_5605(II22745,g14725);
  not NOT_5606(g16733,II22745);
  not NOT_5607(g16739,g14922);
  not NOT_5608(g16743,g14936);
  not NOT_5609(g16749,g15782);
  not NOT_5610(II22752,g14657);
  not NOT_5611(g16758,II22752);
  not NOT_5612(II22755,g14650);
  not NOT_5613(g16761,II22755);
  not NOT_5614(g16764,g14976);
  not NOT_5615(II22759,g14703);
  not NOT_5616(g16767,II22759);
  not NOT_5617(g16770,g14991);
  not NOT_5618(II22763,g14753);
  not NOT_5619(g16775,II22763);
  not NOT_5620(g16781,g15003);
  not NOT_5621(II22768,g14691);
  not NOT_5622(g16785,II22768);
  not NOT_5623(II22771,g14677);
  not NOT_5624(g16788,II22771);
  not NOT_5625(g16791,g15065);
  not NOT_5626(II22775,g14737);
  not NOT_5627(g16794,II22775);
  not NOT_5628(g16797,g15080);
  not NOT_5629(g16804,g15803);
  not NOT_5630(g16809,g15842);
  not NOT_5631(II22783,g13572);
  not NOT_5632(g16813,II22783);
  not NOT_5633(II22786,g14725);
  not NOT_5634(g16814,II22786);
  not NOT_5635(II22789,g14711);
  not NOT_5636(g16817,II22789);
  not NOT_5637(g16820,g15161);
  not NOT_5638(g16825,g15855);
  not NOT_5639(II22797,g14165);
  not NOT_5640(g16830,II22797);
  not NOT_5641(II22800,g13581);
  not NOT_5642(g16831,II22800);
  not NOT_5643(II22803,g14753);
  not NOT_5644(g16832,II22803);
  not NOT_5645(g16836,g15818);
  not NOT_5646(g16840,g15878);
  not NOT_5647(II22810,g14280);
  not NOT_5648(g16842,II22810);
  not NOT_5649(II22813,g13601);
  not NOT_5650(g16843,II22813);
  not NOT_5651(g16846,g15903);
  not NOT_5652(II22820,g14402);
  not NOT_5653(g16848,II22820);
  not NOT_5654(II22823,g13613);
  not NOT_5655(g16849,II22823);
  not NOT_5656(II22828,g14514);
  not NOT_5657(g16852,II22828);
  not NOT_5658(II22836,g13571);
  not NOT_5659(g16858,II22836);
  not NOT_5660(II22842,g13580);
  not NOT_5661(g16862,II22842);
  not NOT_5662(II22845,g13579);
  not NOT_5663(g16863,II22845);
  not NOT_5664(g16867,g13589);
  not NOT_5665(II22852,g13600);
  not NOT_5666(g16877,II22852);
  not NOT_5667(II22855,g13588);
  not NOT_5668(g16878,II22855);
  not NOT_5669(II22860,g14885);
  not NOT_5670(g16881,II22860);
  not NOT_5671(g16884,g13589);
  not NOT_5672(g16895,g13589);
  not NOT_5673(II22866,g13612);
  not NOT_5674(g16905,II22866);
  not NOT_5675(II22869,g13608);
  not NOT_5676(g16906,II22869);
  not NOT_5677(II22875,g14966);
  not NOT_5678(g16910,II22875);
  not NOT_5679(g16913,g13589);
  not NOT_5680(g16924,g13589);
  not NOT_5681(II22881,g13622);
  not NOT_5682(g16934,II22881);
  not NOT_5683(II22893,g15055);
  not NOT_5684(g16940,II22893);
  not NOT_5685(g16943,g13589);
  not NOT_5686(g16954,g13589);
  not NOT_5687(II22912,g15151);
  not NOT_5688(g16971,II22912);
  not NOT_5689(g16974,g13589);
  not NOT_5690(g17029,g14685);
  not NOT_5691(g17057,g13519);
  not NOT_5692(g17063,g14719);
  not NOT_5693(g17092,g13530);
  not NOT_5694(g17098,g14747);
  not NOT_5695(g17130,g13541);
  not NOT_5696(g17136,g14768);
  not NOT_5697(g17157,g13552);
  not NOT_5698(II23253,g13741);
  not NOT_5699(g17189,II23253);
  not NOT_5700(II23274,g13741);
  not NOT_5701(g17200,II23274);
  not NOT_5702(g17203,g13568);
  not NOT_5703(II23287,g13741);
  not NOT_5704(g17207,II23287);
  not NOT_5705(g17208,g13576);
  not NOT_5706(II23292,g13741);
  not NOT_5707(g17212,II23292);
  not NOT_5708(g17214,g13585);
  not NOT_5709(g17217,g13605);
  not NOT_5710(II23309,g16132);
  not NOT_5711(g17227,II23309);
  not NOT_5712(II23314,g15720);
  not NOT_5713(g17230,II23314);
  not NOT_5714(II23317,g16181);
  not NOT_5715(g17233,II23317);
  not NOT_5716(II23323,g15664);
  not NOT_5717(g17237,II23323);
  not NOT_5718(II23326,g15758);
  not NOT_5719(g17240,II23326);
  not NOT_5720(II23329,g15760);
  not NOT_5721(g17243,II23329);
  not NOT_5722(II23335,g16412);
  not NOT_5723(g17249,II23335);
  not NOT_5724(II23338,g15721);
  not NOT_5725(g17252,II23338);
  not NOT_5726(II23341,g15784);
  not NOT_5727(g17255,II23341);
  not NOT_5728(g17258,g16053);
  not NOT_5729(II23345,g15723);
  not NOT_5730(g17259,II23345);
  not NOT_5731(II23348,g15786);
  not NOT_5732(g17262,II23348);
  not NOT_5733(II23351,g15788);
  not NOT_5734(g17265,II23351);
  not NOT_5735(II23358,g16442);
  not NOT_5736(g17272,II23358);
  not NOT_5737(II23361,g15759);
  not NOT_5738(g17275,II23361);
  not NOT_5739(II23364,g15805);
  not NOT_5740(g17278,II23364);
  not NOT_5741(g17281,g16081);
  not NOT_5742(II23368,g16446);
  not NOT_5743(g17282,II23368);
  not NOT_5744(II23371,g15761);
  not NOT_5745(g17285,II23371);
  not NOT_5746(II23374,g15807);
  not NOT_5747(g17288,II23374);
  not NOT_5748(II23377,g15763);
  not NOT_5749(g17291,II23377);
  not NOT_5750(II23380,g15809);
  not NOT_5751(g17294,II23380);
  not NOT_5752(II23383,g15811);
  not NOT_5753(g17297,II23383);
  not NOT_5754(II23386,g13469);
  not NOT_5755(g17300,II23386);
  not NOT_5756(II23392,g13476);
  not NOT_5757(g17304,II23392);
  not NOT_5758(II23395,g15785);
  not NOT_5759(g17307,II23395);
  not NOT_5760(II23398,g15820);
  not NOT_5761(g17310,II23398);
  not NOT_5762(g17313,g16109);
  not NOT_5763(g17314,g16110);
  not NOT_5764(II23403,g13478);
  not NOT_5765(g17315,II23403);
  not NOT_5766(II23406,g15787);
  not NOT_5767(g17318,II23406);
  not NOT_5768(II23409,g15822);
  not NOT_5769(g17321,II23409);
  not NOT_5770(II23412,g13482);
  not NOT_5771(g17324,II23412);
  not NOT_5772(II23415,g15789);
  not NOT_5773(g17327,II23415);
  not NOT_5774(II23418,g15824);
  not NOT_5775(g17330,II23418);
  not NOT_5776(II23421,g15791);
  not NOT_5777(g17333,II23421);
  not NOT_5778(II23424,g15826);
  not NOT_5779(g17336,II23424);
  not NOT_5780(II23430,g13494);
  not NOT_5781(g17342,II23430);
  not NOT_5782(II23433,g15806);
  not NOT_5783(g17345,II23433);
  not NOT_5784(II23436,g15832);
  not NOT_5785(g17348,II23436);
  not NOT_5786(g17351,g16152);
  not NOT_5787(II23442,g13495);
  not NOT_5788(g17354,II23442);
  not NOT_5789(II23445,g15808);
  not NOT_5790(g17357,II23445);
  not NOT_5791(II23448,g15834);
  not NOT_5792(g17360,II23448);
  not NOT_5793(II23451,g13497);
  not NOT_5794(g17363,II23451);
  not NOT_5795(II23454,g15810);
  not NOT_5796(g17366,II23454);
  not NOT_5797(II23457,g15836);
  not NOT_5798(g17369,II23457);
  not NOT_5799(II23460,g13501);
  not NOT_5800(g17372,II23460);
  not NOT_5801(II23463,g15812);
  not NOT_5802(g17375,II23463);
  not NOT_5803(II23466,g15838);
  not NOT_5804(g17378,II23466);
  not NOT_5805(II23472,g13510);
  not NOT_5806(g17384,II23472);
  not NOT_5807(II23475,g15821);
  not NOT_5808(g17387,II23475);
  not NOT_5809(II23478,g15844);
  not NOT_5810(g17390,II23478);
  not NOT_5811(g17394,g16197);
  not NOT_5812(II23487,g13511);
  not NOT_5813(g17399,II23487);
  not NOT_5814(II23490,g15823);
  not NOT_5815(g17402,II23490);
  not NOT_5816(II23493,g15846);
  not NOT_5817(g17405,II23493);
  not NOT_5818(II23498,g13512);
  not NOT_5819(g17410,II23498);
  not NOT_5820(II23501,g15825);
  not NOT_5821(g17413,II23501);
  not NOT_5822(II23504,g15848);
  not NOT_5823(g17416,II23504);
  not NOT_5824(II23507,g13514);
  not NOT_5825(g17419,II23507);
  not NOT_5826(II23510,g15827);
  not NOT_5827(g17422,II23510);
  not NOT_5828(II23513,g15850);
  not NOT_5829(g17425,II23513);
  not NOT_5830(II23518,g15856);
  not NOT_5831(g17430,II23518);
  not NOT_5832(II23521,g13518);
  not NOT_5833(g17433,II23521);
  not NOT_5834(II23524,g15833);
  not NOT_5835(g17436,II23524);
  not NOT_5836(II23527,g15858);
  not NOT_5837(g17439,II23527);
  not NOT_5838(II23530,g14885);
  not NOT_5839(g17442,II23530);
  not NOT_5840(g17445,g16250);
  not NOT_5841(II23539,g13524);
  not NOT_5842(g17451,II23539);
  not NOT_5843(II23542,g15835);
  not NOT_5844(g17454,II23542);
  not NOT_5845(II23545,g15867);
  not NOT_5846(g17457,II23545);
  not NOT_5847(II23553,g13525);
  not NOT_5848(g17465,II23553);
  not NOT_5849(II23556,g15837);
  not NOT_5850(g17468,II23556);
  not NOT_5851(II23559,g15869);
  not NOT_5852(g17471,II23559);
  not NOT_5853(II23564,g13526);
  not NOT_5854(g17476,II23564);
  not NOT_5855(II23567,g15839);
  not NOT_5856(g17479,II23567);
  not NOT_5857(II23570,g15871);
  not NOT_5858(g17482,II23570);
  not NOT_5859(II23575,g15843);
  not NOT_5860(g17487,II23575);
  not NOT_5861(II23578,g15879);
  not NOT_5862(g17490,II23578);
  not NOT_5863(II23581,g13528);
  not NOT_5864(g17493,II23581);
  not NOT_5865(II23584,g15845);
  not NOT_5866(g17496,II23584);
  not NOT_5867(g17499,g16292);
  not NOT_5868(II23588,g14885);
  not NOT_5869(g17500,II23588);
  not NOT_5870(II23591,g14885);
  not NOT_5871(g17503,II23591);
  not NOT_5872(II23599,g15887);
  not NOT_5873(g17511,II23599);
  not NOT_5874(II23602,g13529);
  not NOT_5875(g17514,II23602);
  not NOT_5876(II23605,g15847);
  not NOT_5877(g17517,II23605);
  not NOT_5878(II23608,g15889);
  not NOT_5879(g17520,II23608);
  not NOT_5880(II23611,g14966);
  not NOT_5881(g17523,II23611);
  not NOT_5882(II23619,g13535);
  not NOT_5883(g17531,II23619);
  not NOT_5884(II23622,g15849);
  not NOT_5885(g17534,II23622);
  not NOT_5886(II23625,g15898);
  not NOT_5887(g17537,II23625);
  not NOT_5888(II23633,g13536);
  not NOT_5889(g17545,II23633);
  not NOT_5890(II23636,g15851);
  not NOT_5891(g17548,II23636);
  not NOT_5892(II23639,g15900);
  not NOT_5893(g17551,II23639);
  not NOT_5894(II23645,g13537);
  not NOT_5895(g17557,II23645);
  not NOT_5896(II23648,g15857);
  not NOT_5897(g17560,II23648);
  not NOT_5898(II23651,g13538);
  not NOT_5899(g17563,II23651);
  not NOT_5900(g17566,g16346);
  not NOT_5901(II23655,g14831);
  not NOT_5902(g17567,II23655);
  not NOT_5903(II23658,g14885);
  not NOT_5904(g17570,II23658);
  not NOT_5905(II23661,g16085);
  not NOT_5906(g17573,II23661);
  not NOT_5907(II23667,g15866);
  not NOT_5908(g17579,II23667);
  not NOT_5909(II23670,g15912);
  not NOT_5910(g17582,II23670);
  not NOT_5911(II23673,g13539);
  not NOT_5912(g17585,II23673);
  not NOT_5913(II23676,g15868);
  not NOT_5914(g17588,II23676);
  not NOT_5915(II23679,g14966);
  not NOT_5916(g17591,II23679);
  not NOT_5917(II23682,g14966);
  not NOT_5918(g17594,II23682);
  not NOT_5919(II23689,g15920);
  not NOT_5920(g17601,II23689);
  not NOT_5921(II23692,g13540);
  not NOT_5922(g17604,II23692);
  not NOT_5923(II23695,g15870);
  not NOT_5924(g17607,II23695);
  not NOT_5925(II23698,g15922);
  not NOT_5926(g17610,II23698);
  not NOT_5927(II23701,g15055);
  not NOT_5928(g17613,II23701);
  not NOT_5929(II23709,g13546);
  not NOT_5930(g17621,II23709);
  not NOT_5931(II23712,g15872);
  not NOT_5932(g17624,II23712);
  not NOT_5933(II23715,g15931);
  not NOT_5934(g17627,II23715);
  not NOT_5935(II23725,g13547);
  not NOT_5936(g17637,II23725);
  not NOT_5937(g17640,g13873);
  not NOT_5938(II23729,g14337);
  not NOT_5939(g17645,II23729);
  not NOT_5940(g17648,g16384);
  not NOT_5941(II23733,g14831);
  not NOT_5942(g17649,II23733);
  not NOT_5943(II23739,g13548);
  not NOT_5944(g17655,II23739);
  not NOT_5945(II23742,g15888);
  not NOT_5946(g17658,II23742);
  not NOT_5947(II23745,g13549);
  not NOT_5948(g17661,II23745);
  not NOT_5949(II23748,g14904);
  not NOT_5950(g17664,II23748);
  not NOT_5951(II23751,g14966);
  not NOT_5952(g17667,II23751);
  not NOT_5953(II23754,g16123);
  not NOT_5954(g17670,II23754);
  not NOT_5955(II23760,g15897);
  not NOT_5956(g17676,II23760);
  not NOT_5957(II23763,g15941);
  not NOT_5958(g17679,II23763);
  not NOT_5959(II23766,g13550);
  not NOT_5960(g17682,II23766);
  not NOT_5961(II23769,g15899);
  not NOT_5962(g17685,II23769);
  not NOT_5963(II23772,g15055);
  not NOT_5964(g17688,II23772);
  not NOT_5965(II23775,g15055);
  not NOT_5966(g17691,II23775);
  not NOT_5967(II23782,g15949);
  not NOT_5968(g17698,II23782);
  not NOT_5969(II23785,g13551);
  not NOT_5970(g17701,II23785);
  not NOT_5971(II23788,g15901);
  not NOT_5972(g17704,II23788);
  not NOT_5973(II23791,g15951);
  not NOT_5974(g17707,II23791);
  not NOT_5975(II23794,g15151);
  not NOT_5976(g17710,II23794);
  not NOT_5977(g17720,g15853);
  not NOT_5978(g17724,g13886);
  not NOT_5979(II23817,g13557);
  not NOT_5980(g17738,II23817);
  not NOT_5981(g17741,g13895);
  not NOT_5982(II23821,g14337);
  not NOT_5983(g17746,II23821);
  not NOT_5984(II23824,g14904);
  not NOT_5985(g17749,II23824);
  not NOT_5986(II23830,g13558);
  not NOT_5987(g17755,II23830);
  not NOT_5988(II23833,g15921);
  not NOT_5989(g17758,II23833);
  not NOT_5990(II23836,g13559);
  not NOT_5991(g17761,II23836);
  not NOT_5992(II23839,g14985);
  not NOT_5993(g17764,II23839);
  not NOT_5994(II23842,g15055);
  not NOT_5995(g17767,II23842);
  not NOT_5996(II23845,g16174);
  not NOT_5997(g17770,II23845);
  not NOT_5998(II23851,g15930);
  not NOT_5999(g17776,II23851);
  not NOT_6000(II23854,g15970);
  not NOT_6001(g17779,II23854);
  not NOT_6002(II23857,g13560);
  not NOT_6003(g17782,II23857);
  not NOT_6004(II23860,g15932);
  not NOT_6005(g17785,II23860);
  not NOT_6006(II23863,g15151);
  not NOT_6007(g17788,II23863);
  not NOT_6008(II23866,g15151);
  not NOT_6009(g17791,II23866);
  not NOT_6010(II23874,g15797);
  not NOT_6011(g17799,II23874);
  not NOT_6012(g17802,g13907);
  not NOT_6013(II23888,g14685);
  not NOT_6014(g17815,II23888);
  not NOT_6015(g17825,g13927);
  not NOT_6016(II23904,g13561);
  not NOT_6017(g17839,II23904);
  not NOT_6018(g17842,g13936);
  not NOT_6019(II23908,g14337);
  not NOT_6020(g17847,II23908);
  not NOT_6021(II23911,g14985);
  not NOT_6022(g17850,II23911);
  not NOT_6023(II23917,g13562);
  not NOT_6024(g17856,II23917);
  not NOT_6025(II23920,g15950);
  not NOT_6026(g17859,II23920);
  not NOT_6027(II23923,g13563);
  not NOT_6028(g17862,II23923);
  not NOT_6029(II23926,g15074);
  not NOT_6030(g17865,II23926);
  not NOT_6031(II23929,g15151);
  not NOT_6032(g17868,II23929);
  not NOT_6033(II23932,g16233);
  not NOT_6034(g17871,II23932);
  not NOT_6035(g17878,g15830);
  not NOT_6036(g17882,g13946);
  not NOT_6037(g17892,g13954);
  not NOT_6038(g17893,g14165);
  not NOT_6039(II23954,g16154);
  not NOT_6040(g17903,II23954);
  not NOT_6041(g17914,g13963);
  not NOT_6042(II23976,g14719);
  not NOT_6043(g17927,II23976);
  not NOT_6044(g17937,g13983);
  not NOT_6045(II23992,g13564);
  not NOT_6046(g17951,II23992);
  not NOT_6047(g17954,g13992);
  not NOT_6048(II23996,g14337);
  not NOT_6049(g17959,II23996);
  not NOT_6050(II23999,g15074);
  not NOT_6051(g17962,II23999);
  not NOT_6052(g17969,g15841);
  not NOT_6053(g17974,g14001);
  not NOT_6054(g17984,g14008);
  not NOT_6055(g17988,g14685);
  not NOT_6056(g17991,g14450);
  not NOT_6057(g17993,g14016);
  not NOT_6058(g18003,g14024);
  not NOT_6059(g18004,g14280);
  not NOT_6060(II24049,g16213);
  not NOT_6061(g18014,II24049);
  not NOT_6062(g18025,g14033);
  not NOT_6063(II24071,g14747);
  not NOT_6064(g18038,II24071);
  not NOT_6065(g18048,g14053);
  not NOT_6066(g18063,g15660);
  not NOT_6067(g18070,g15854);
  not NOT_6068(g18074,g14062);
  not NOT_6069(g18084,g14068);
  not NOT_6070(g18089,g14355);
  not NOT_6071(g18091,g14092);
  not NOT_6072(g18101,g14099);
  not NOT_6073(g18105,g14719);
  not NOT_6074(g18108,g14537);
  not NOT_6075(g18110,g14107);
  not NOT_6076(g18120,g14115);
  not NOT_6077(g18121,g14402);
  not NOT_6078(II24144,g16278);
  not NOT_6079(g18131,II24144);
  not NOT_6080(g18142,g14124);
  not NOT_6081(II24166,g14768);
  not NOT_6082(g18155,II24166);
  not NOT_6083(II24171,g16439);
  not NOT_6084(g18166,II24171);
  not NOT_6085(g18170,g15877);
  not NOT_6086(g18174,g14148);
  not NOT_6087(g18179,g14153);
  not NOT_6088(g18188,g14252);
  not NOT_6089(g18190,g14177);
  not NOT_6090(g18200,g14183);
  not NOT_6091(g18205,g14467);
  not NOT_6092(g18207,g14207);
  not NOT_6093(g18217,g14214);
  not NOT_6094(g18221,g14747);
  not NOT_6095(g18224,g14592);
  not NOT_6096(g18226,g14222);
  not NOT_6097(g18236,g14230);
  not NOT_6098(g18237,g14514);
  not NOT_6099(II24247,g16337);
  not NOT_6100(g18247,II24247);
  not NOT_6101(II24258,g16463);
  not NOT_6102(g18258,II24258);
  not NOT_6103(g18261,g15719);
  not NOT_6104(g18265,g14238);
  not NOT_6105(g18275,g14171);
  not NOT_6106(II24285,g15992);
  not NOT_6107(g18278,II24285);
  not NOT_6108(g18281,g14263);
  not NOT_6109(g18286,g14268);
  not NOT_6110(g18295,g14374);
  not NOT_6111(g18297,g14292);
  not NOT_6112(g18307,g14298);
  not NOT_6113(g18312,g14554);
  not NOT_6114(g18314,g14322);
  not NOT_6115(g18324,g14329);
  not NOT_6116(g18328,g14768);
  not NOT_6117(g18331,g14626);
  not NOT_6118(II24346,g15873);
  not NOT_6119(g18334,II24346);
  not NOT_6120(g18337,g15757);
  not NOT_6121(g18341,g14342);
  not NOT_6122(g18351,g13741);
  not NOT_6123(g18353,g13918);
  not NOT_6124(II24368,g15990);
  not NOT_6125(g18355,II24368);
  not NOT_6126(g18358,g14360);
  not NOT_6127(g18368,g14286);
  not NOT_6128(II24394,g15995);
  not NOT_6129(g18371,II24394);
  not NOT_6130(g18374,g14385);
  not NOT_6131(g18379,g14390);
  not NOT_6132(g18388,g14486);
  not NOT_6133(g18390,g14414);
  not NOT_6134(g18400,g14420);
  not NOT_6135(g18405,g14609);
  not NOT_6136(g18407,g15959);
  not NOT_6137(g18414,g15718);
  not NOT_6138(g18415,g15783);
  not NOT_6139(g18429,g14831);
  not NOT_6140(II24459,g13599);
  not NOT_6141(g18432,II24459);
  not NOT_6142(g18435,g14359);
  not NOT_6143(g18436,g14454);
  not NOT_6144(g18446,g13741);
  not NOT_6145(g18448,g13974);
  not NOT_6146(II24481,g15993);
  not NOT_6147(g18450,II24481);
  not NOT_6148(g18453,g14472);
  not NOT_6149(g18463,g14408);
  not NOT_6150(II24507,g15999);
  not NOT_6151(g18466,II24507);
  not NOT_6152(g18469,g14497);
  not NOT_6153(g18474,g14502);
  not NOT_6154(g18483,g14573);
  not NOT_6155(g18485,g15756);
  not NOT_6156(g18486,g15804);
  not NOT_6157(g18490,g13565);
  not NOT_6158(g18502,g14904);
  not NOT_6159(II24560,g13611);
  not NOT_6160(g18505,II24560);
  not NOT_6161(g18508,g14471);
  not NOT_6162(g18509,g14541);
  not NOT_6163(g18519,g13741);
  not NOT_6164(g18521,g14044);
  not NOT_6165(II24582,g15996);
  not NOT_6166(g18523,II24582);
  not NOT_6167(g18526,g14559);
  not NOT_6168(g18536,g14520);
  not NOT_6169(II24608,g16006);
  not NOT_6170(g18539,II24608);
  not NOT_6171(g18543,g15819);
  not NOT_6172(g18552,g16154);
  not NOT_6173(g18554,g13573);
  not NOT_6174(g18566,g14985);
  not NOT_6175(II24662,g13621);
  not NOT_6176(g18569,II24662);
  not NOT_6177(g18572,g14558);
  not NOT_6178(g18573,g14596);
  not NOT_6179(g18583,g13741);
  not NOT_6180(g18585,g14135);
  not NOT_6181(II24684,g16000);
  not NOT_6182(g18587,II24684);
  not NOT_6183(g18593,g15831);
  not NOT_6184(g18602,g16213);
  not NOT_6185(g18604,g13582);
  not NOT_6186(g18616,g15074);
  not NOT_6187(II24732,g13633);
  not NOT_6188(g18619,II24732);
  not NOT_6189(g18622,g14613);
  not NOT_6190(g18634,g16278);
  not NOT_6191(g18636,g13602);
  not NOT_6192(g18643,g16337);
  not NOT_6193(g18646,g16341);
  not NOT_6194(g18656,g14776);
  not NOT_6195(g18670,g14797);
  not NOT_6196(g18679,g14811);
  not NOT_6197(g18691,g14885);
  not NOT_6198(g18692,g14837);
  not NOT_6199(g18699,g14849);
  not NOT_6200(g18708,g14863);
  not NOT_6201(g18720,g14895);
  not NOT_6202(g18725,g13865);
  not NOT_6203(g18727,g14966);
  not NOT_6204(g18728,g14910);
  not NOT_6205(g18735,g14922);
  not NOT_6206(g18744,g14936);
  not NOT_6207(g18756,g14960);
  not NOT_6208(g18757,g14963);
  not NOT_6209(g18758,g14976);
  not NOT_6210(g18764,g15055);
  not NOT_6211(g18765,g14991);
  not NOT_6212(g18772,g15003);
  not NOT_6213(g18783,g15034);
  not NOT_6214(g18784,g15037);
  not NOT_6215(g18785,g15040);
  not NOT_6216(g18786,g15043);
  not NOT_6217(g18787,g15049);
  not NOT_6218(g18788,g15052);
  not NOT_6219(g18789,g15065);
  not NOT_6220(g18795,g15151);
  not NOT_6221(g18796,g15080);
  not NOT_6222(g18805,g15106);
  not NOT_6223(g18806,g15109);
  not NOT_6224(g18807,g15112);
  not NOT_6225(g18808,g15115);
  not NOT_6226(g18809,g15130);
  not NOT_6227(g18810,g15133);
  not NOT_6228(g18811,g15136);
  not NOT_6229(g18812,g15139);
  not NOT_6230(g18813,g15145);
  not NOT_6231(g18814,g15148);
  not NOT_6232(g18815,g15161);
  not NOT_6233(g18822,g15179);
  not NOT_6234(g18823,g15182);
  not NOT_6235(g18824,g15185);
  not NOT_6236(g18825,g15198);
  not NOT_6237(g18826,g15201);
  not NOT_6238(g18827,g15204);
  not NOT_6239(g18828,g15207);
  not NOT_6240(g18829,g15222);
  not NOT_6241(g18830,g15225);
  not NOT_6242(g18831,g15228);
  not NOT_6243(g18832,g15231);
  not NOT_6244(g18833,g15237);
  not NOT_6245(g18834,g15240);
  not NOT_6246(g18838,g15248);
  not NOT_6247(g18839,g15251);
  not NOT_6248(g18840,g15254);
  not NOT_6249(g18841,g15265);
  not NOT_6250(g18842,g15268);
  not NOT_6251(g18843,g15271);
  not NOT_6252(g18844,g15284);
  not NOT_6253(g18845,g15287);
  not NOT_6254(g18846,g15290);
  not NOT_6255(g18847,g15293);
  not NOT_6256(g18848,g15308);
  not NOT_6257(g18849,g15311);
  not NOT_6258(g18850,g15314);
  not NOT_6259(g18851,g15317);
  not NOT_6260(g18853,g15326);
  not NOT_6261(g18854,g15329);
  not NOT_6262(g18855,g15332);
  not NOT_6263(g18856,g15340);
  not NOT_6264(g18857,g15343);
  not NOT_6265(g18858,g15346);
  not NOT_6266(g18859,g15357);
  not NOT_6267(g18860,g15360);
  not NOT_6268(g18861,g15363);
  not NOT_6269(g18862,g15376);
  not NOT_6270(g18863,g15379);
  not NOT_6271(g18864,g15382);
  not NOT_6272(g18865,g15385);
  not NOT_6273(II24894,g14797);
  not NOT_6274(g18869,II24894);
  not NOT_6275(g18870,g15393);
  not NOT_6276(g18871,g15396);
  not NOT_6277(g18872,g15399);
  not NOT_6278(g18873,g15404);
  not NOT_6279(g18874,g15412);
  not NOT_6280(g18875,g15415);
  not NOT_6281(g18876,g15418);
  not NOT_6282(g18877,g15426);
  not NOT_6283(g18878,g15429);
  not NOT_6284(g18879,g15432);
  not NOT_6285(g18880,g15443);
  not NOT_6286(g18881,g15446);
  not NOT_6287(g18882,g15449);
  not NOT_6288(g18884,g13469);
  not NOT_6289(II24913,g15800);
  not NOT_6290(g18886,II24913);
  not NOT_6291(II24916,g14776);
  not NOT_6292(g18890,II24916);
  not NOT_6293(g18891,g15461);
  not NOT_6294(g18892,g15464);
  not NOT_6295(g18893,g15467);
  not NOT_6296(g18894,g15471);
  not NOT_6297(II24923,g14849);
  not NOT_6298(g18895,II24923);
  not NOT_6299(g18896,g15477);
  not NOT_6300(g18897,g15480);
  not NOT_6301(g18898,g15483);
  not NOT_6302(g18899,g15488);
  not NOT_6303(g18900,g15496);
  not NOT_6304(g18901,g15499);
  not NOT_6305(g18902,g15502);
  not NOT_6306(g18903,g15510);
  not NOT_6307(g18904,g15513);
  not NOT_6308(g18905,g15516);
  not NOT_6309(g18908,g15521);
  not NOT_6310(g18909,g15528);
  not NOT_6311(g18910,g15531);
  not NOT_6312(g18911,g15534);
  not NOT_6313(g18912,g15537);
  not NOT_6314(II24943,g14811);
  not NOT_6315(g18913,II24943);
  not NOT_6316(g18914,g15547);
  not NOT_6317(g18915,g15550);
  not NOT_6318(g18916,g15553);
  not NOT_6319(g18917,g15557);
  not NOT_6320(II24950,g14922);
  not NOT_6321(g18918,II24950);
  not NOT_6322(g18919,g15563);
  not NOT_6323(g18920,g15566);
  not NOT_6324(g18921,g15569);
  not NOT_6325(g18922,g15574);
  not NOT_6326(g18923,g15582);
  not NOT_6327(g18924,g15585);
  not NOT_6328(g18925,g15588);
  not NOT_6329(g18926,g15596);
  not NOT_6330(g18927,g15599);
  not NOT_6331(g18928,g15606);
  not NOT_6332(g18929,g15609);
  not NOT_6333(g18930,g15612);
  not NOT_6334(g18931,g15615);
  not NOT_6335(II24966,g14863);
  not NOT_6336(g18932,II24966);
  not NOT_6337(g18933,g15625);
  not NOT_6338(g18934,g15628);
  not NOT_6339(g18935,g15631);
  not NOT_6340(g18936,g15635);
  not NOT_6341(II24973,g15003);
  not NOT_6342(g18937,II24973);
  not NOT_6343(g18938,g15641);
  not NOT_6344(g18939,g15644);
  not NOT_6345(g18940,g15647);
  not NOT_6346(g18941,g15652);
  not NOT_6347(g18943,g15655);
  not NOT_6348(II24982,g14347);
  not NOT_6349(g18944,II24982);
  not NOT_6350(g18945,g15667);
  not NOT_6351(g18946,g15672);
  not NOT_6352(g18947,g15675);
  not NOT_6353(g18948,g15682);
  not NOT_6354(g18949,g15685);
  not NOT_6355(g18950,g15688);
  not NOT_6356(g18951,g15691);
  not NOT_6357(II24992,g14936);
  not NOT_6358(g18952,II24992);
  not NOT_6359(g18953,g15701);
  not NOT_6360(g18954,g15704);
  not NOT_6361(g18955,g15707);
  not NOT_6362(g18956,g15711);
  not NOT_6363(g18958,g15714);
  not NOT_6364(II25001,g14244);
  not NOT_6365(g18959,II25001);
  not NOT_6366(II25004,g14459);
  not NOT_6367(g18960,II25004);
  not NOT_6368(g18961,g15726);
  not NOT_6369(g18962,g15731);
  not NOT_6370(g18963,g15734);
  not NOT_6371(g18964,g15741);
  not NOT_6372(g18965,g15744);
  not NOT_6373(g18966,g15747);
  not NOT_6374(g18967,g15750);
  not NOT_6375(II25015,g14158);
  not NOT_6376(g18969,II25015);
  not NOT_6377(II25018,g14366);
  not NOT_6378(g18970,II25018);
  not NOT_6379(II25021,g14546);
  not NOT_6380(g18971,II25021);
  not NOT_6381(g18972,g15766);
  not NOT_6382(g18973,g15771);
  not NOT_6383(g18974,g15774);
  not NOT_6384(g18976,g15777);
  not NOT_6385(II25037,g14071);
  not NOT_6386(g18981,II25037);
  not NOT_6387(II25041,g14895);
  not NOT_6388(g18983,II25041);
  not NOT_6389(II25044,g14273);
  not NOT_6390(g18984,II25044);
  not NOT_6391(II25047,g14478);
  not NOT_6392(g18985,II25047);
  not NOT_6393(II25050,g14601);
  not NOT_6394(g18986,II25050);
  not NOT_6395(g18987,g15794);
  not NOT_6396(II25054,g14837);
  not NOT_6397(g18988,II25054);
  not NOT_6398(II25057,g14186);
  not NOT_6399(g18989,II25057);
  not NOT_6400(II25061,g14976);
  not NOT_6401(g18991,II25061);
  not NOT_6402(II25064,g14395);
  not NOT_6403(g18992,II25064);
  not NOT_6404(II25067,g14565);
  not NOT_6405(g18993,II25067);
  not NOT_6406(II25071,g14910);
  not NOT_6407(g18995,II25071);
  not NOT_6408(II25074,g14301);
  not NOT_6409(g18996,II25074);
  not NOT_6410(II25078,g15065);
  not NOT_6411(g18998,II25078);
  not NOT_6412(II25081,g14507);
  not NOT_6413(g18999,II25081);
  not NOT_6414(II25084,g14885);
  not NOT_6415(g19000,II25084);
  not NOT_6416(g19001,g14071);
  not NOT_6417(II25089,g14991);
  not NOT_6418(g19008,II25089);
  not NOT_6419(II25092,g14423);
  not NOT_6420(g19009,II25092);
  not NOT_6421(II25096,g15161);
  not NOT_6422(g19011,II25096);
  not NOT_6423(II25099,g19000);
  not NOT_6424(g19012,II25099);
  not NOT_6425(II25102,g18944);
  not NOT_6426(g19013,II25102);
  not NOT_6427(II25105,g18959);
  not NOT_6428(g19014,II25105);
  not NOT_6429(II25108,g18969);
  not NOT_6430(g19015,II25108);
  not NOT_6431(II25111,g18981);
  not NOT_6432(g19016,II25111);
  not NOT_6433(II25114,g18983);
  not NOT_6434(g19017,II25114);
  not NOT_6435(II25117,g18988);
  not NOT_6436(g19018,II25117);
  not NOT_6437(II25120,g18869);
  not NOT_6438(g19019,II25120);
  not NOT_6439(II25123,g18890);
  not NOT_6440(g19020,II25123);
  not NOT_6441(II25126,g16858);
  not NOT_6442(g19021,II25126);
  not NOT_6443(II25129,g16813);
  not NOT_6444(g19022,II25129);
  not NOT_6445(II25132,g16862);
  not NOT_6446(g19023,II25132);
  not NOT_6447(II25135,g16506);
  not NOT_6448(g19024,II25135);
  not NOT_6449(II25138,g18960);
  not NOT_6450(g19025,II25138);
  not NOT_6451(II25141,g18970);
  not NOT_6452(g19026,II25141);
  not NOT_6453(II25144,g18984);
  not NOT_6454(g19027,II25144);
  not NOT_6455(II25147,g18989);
  not NOT_6456(g19028,II25147);
  not NOT_6457(II25150,g18991);
  not NOT_6458(g19029,II25150);
  not NOT_6459(II25153,g18995);
  not NOT_6460(g19030,II25153);
  not NOT_6461(II25156,g18895);
  not NOT_6462(g19031,II25156);
  not NOT_6463(II25159,g18913);
  not NOT_6464(g19032,II25159);
  not NOT_6465(II25162,g16863);
  not NOT_6466(g19033,II25162);
  not NOT_6467(II25165,g16831);
  not NOT_6468(g19034,II25165);
  not NOT_6469(II25168,g16877);
  not NOT_6470(g19035,II25168);
  not NOT_6471(II25171,g16528);
  not NOT_6472(g19036,II25171);
  not NOT_6473(II25174,g18971);
  not NOT_6474(g19037,II25174);
  not NOT_6475(II25177,g18985);
  not NOT_6476(g19038,II25177);
  not NOT_6477(II25180,g18992);
  not NOT_6478(g19039,II25180);
  not NOT_6479(II25183,g18996);
  not NOT_6480(g19040,II25183);
  not NOT_6481(II25186,g18998);
  not NOT_6482(g19041,II25186);
  not NOT_6483(II25189,g19008);
  not NOT_6484(g19042,II25189);
  not NOT_6485(II25192,g18918);
  not NOT_6486(g19043,II25192);
  not NOT_6487(II25195,g18932);
  not NOT_6488(g19044,II25195);
  not NOT_6489(II25198,g16878);
  not NOT_6490(g19045,II25198);
  not NOT_6491(II25201,g16843);
  not NOT_6492(g19046,II25201);
  not NOT_6493(II25204,g16905);
  not NOT_6494(g19047,II25204);
  not NOT_6495(II25207,g16559);
  not NOT_6496(g19048,II25207);
  not NOT_6497(II25210,g18986);
  not NOT_6498(g19049,II25210);
  not NOT_6499(II25213,g18993);
  not NOT_6500(g19050,II25213);
  not NOT_6501(II25216,g18999);
  not NOT_6502(g19051,II25216);
  not NOT_6503(II25219,g19009);
  not NOT_6504(g19052,II25219);
  not NOT_6505(II25222,g19011);
  not NOT_6506(g19053,II25222);
  not NOT_6507(II25225,g16514);
  not NOT_6508(g19054,II25225);
  not NOT_6509(II25228,g18937);
  not NOT_6510(g19055,II25228);
  not NOT_6511(II25231,g18952);
  not NOT_6512(g19056,II25231);
  not NOT_6513(II25234,g16906);
  not NOT_6514(g19057,II25234);
  not NOT_6515(II25237,g16849);
  not NOT_6516(g19058,II25237);
  not NOT_6517(II25240,g16934);
  not NOT_6518(g19059,II25240);
  not NOT_6519(II25243,g17227);
  not NOT_6520(g19060,II25243);
  not NOT_6521(II25246,g17233);
  not NOT_6522(g19061,II25246);
  not NOT_6523(II25249,g17300);
  not NOT_6524(g19062,II25249);
  not NOT_6525(II25253,g17124);
  not NOT_6526(g19064,II25253);
  not NOT_6527(g19070,g18583);
  not NOT_6528(II25258,g16974);
  not NOT_6529(g19075,II25258);
  not NOT_6530(g19078,g18619);
  not NOT_6531(II25264,g17151);
  not NOT_6532(g19081,II25264);
  not NOT_6533(II25272,g17051);
  not NOT_6534(g19091,II25272);
  not NOT_6535(g19096,g18980);
  not NOT_6536(II25283,g17086);
  not NOT_6537(g19098,II25283);
  not NOT_6538(II25294,g17124);
  not NOT_6539(g19105,II25294);
  not NOT_6540(II25303,g17151);
  not NOT_6541(g19110,II25303);
  not NOT_6542(II25308,g16867);
  not NOT_6543(g19113,II25308);
  not NOT_6544(II25315,g16895);
  not NOT_6545(g19118,II25315);
  not NOT_6546(II25320,g16924);
  not NOT_6547(g19125,II25320);
  not NOT_6548(II25325,g16954);
  not NOT_6549(g19132,II25325);
  not NOT_6550(II25334,g17645);
  not NOT_6551(g19145,II25334);
  not NOT_6552(II25338,g17746);
  not NOT_6553(g19147,II25338);
  not NOT_6554(II25344,g17847);
  not NOT_6555(g19151,II25344);
  not NOT_6556(II25351,g17959);
  not NOT_6557(g19156,II25351);
  not NOT_6558(II25355,g18669);
  not NOT_6559(g19158,II25355);
  not NOT_6560(II25358,g18678);
  not NOT_6561(g19159,II25358);
  not NOT_6562(II25365,g18707);
  not NOT_6563(g19164,II25365);
  not NOT_6564(II25371,g18719);
  not NOT_6565(g19168,II25371);
  not NOT_6566(II25374,g18726);
  not NOT_6567(g19169,II25374);
  not NOT_6568(II25377,g18743);
  not NOT_6569(g19170,II25377);
  not NOT_6570(II25383,g18755);
  not NOT_6571(g19174,II25383);
  not NOT_6572(II25386,g18763);
  not NOT_6573(g19175,II25386);
  not NOT_6574(II25389,g18780);
  not NOT_6575(g19176,II25389);
  not NOT_6576(II25395,g18782);
  not NOT_6577(g19180,II25395);
  not NOT_6578(II25399,g18794);
  not NOT_6579(g19182,II25399);
  not NOT_6580(II25402,g18821);
  not NOT_6581(g19183,II25402);
  not NOT_6582(II25406,g18804);
  not NOT_6583(g19185,II25406);
  not NOT_6584(II25412,g18820);
  not NOT_6585(g19189,II25412);
  not NOT_6586(II25415,g18835);
  not NOT_6587(g19190,II25415);
  not NOT_6588(II25423,g18852);
  not NOT_6589(g19196,II25423);
  not NOT_6590(II25426,g18836);
  not NOT_6591(g19197,II25426);
  not NOT_6592(II25429,g18975);
  not NOT_6593(g19198,II25429);
  not NOT_6594(II25432,g18837);
  not NOT_6595(g19199,II25432);
  not NOT_6596(II25442,g18866);
  not NOT_6597(g19207,II25442);
  not NOT_6598(II25445,g18968);
  not NOT_6599(g19208,II25445);
  not NOT_6600(II25456,g18883);
  not NOT_6601(g19217,II25456);
  not NOT_6602(II25459,g18867);
  not NOT_6603(g19218,II25459);
  not NOT_6604(II25463,g18868);
  not NOT_6605(g19220,II25463);
  not NOT_6606(II25474,g18885);
  not NOT_6607(g19229,II25474);
  not NOT_6608(II25486,g18754);
  not NOT_6609(g19237,II25486);
  not NOT_6610(II25489,g18906);
  not NOT_6611(g19238,II25489);
  not NOT_6612(II25492,g18907);
  not NOT_6613(g19239,II25492);
  not NOT_6614(II25506,g18781);
  not NOT_6615(g19247,II25506);
  not NOT_6616(II25510,g18542);
  not NOT_6617(g19249,II25510);
  not NOT_6618(g19251,g16540);
  not NOT_6619(II25525,g18803);
  not NOT_6620(g19258,II25525);
  not NOT_6621(II25528,g18942);
  not NOT_6622(g19259,II25528);
  not NOT_6623(g19265,g16572);
  not NOT_6624(II25557,g18957);
  not NOT_6625(g19270,II25557);
  not NOT_6626(II25567,g17186);
  not NOT_6627(g19272,II25567);
  not NOT_6628(g19280,g16596);
  not NOT_6629(g19287,g16608);
  not NOT_6630(II25612,g17197);
  not NOT_6631(g19291,II25612);
  not NOT_6632(g19299,g16616);
  not NOT_6633(g19301,g16622);
  not NOT_6634(g19302,g17025);
  not NOT_6635(g19305,g16626);
  not NOT_6636(II25660,g17204);
  not NOT_6637(g19309,II25660);
  not NOT_6638(g19319,g16633);
  not NOT_6639(g19322,g16636);
  not NOT_6640(g19323,g17059);
  not NOT_6641(g19326,g16640);
  not NOT_6642(II25717,g17209);
  not NOT_6643(g19330,II25717);
  not NOT_6644(II25728,g17118);
  not NOT_6645(g19335,II25728);
  not NOT_6646(g19346,g16644);
  not NOT_6647(g19349,g16647);
  not NOT_6648(g19350,g17094);
  not NOT_6649(g19353,g16651);
  not NOT_6650(II25768,g17139);
  not NOT_6651(g19358,II25768);
  not NOT_6652(II25778,g17145);
  not NOT_6653(g19369,II25778);
  not NOT_6654(g19380,g16656);
  not NOT_6655(g19383,g16659);
  not NOT_6656(g19384,g17132);
  not NOT_6657(g19387,g16567);
  not NOT_6658(g19388,g17139);
  not NOT_6659(II25816,g17162);
  not NOT_6660(g19390,II25816);
  not NOT_6661(II25826,g17168);
  not NOT_6662(g19401,II25826);
  not NOT_6663(g19412,g16673);
  not NOT_6664(g19415,g16676);
  not NOT_6665(g19417,g16591);
  not NOT_6666(g19418,g17162);
  not NOT_6667(II25862,g17177);
  not NOT_6668(g19420,II25862);
  not NOT_6669(II25872,g17183);
  not NOT_6670(g19431,II25872);
  not NOT_6671(g19441,g17213);
  not NOT_6672(g19444,g17985);
  not NOT_6673(g19448,g16694);
  not NOT_6674(g19452,g16702);
  not NOT_6675(g19454,g16611);
  not NOT_6676(g19455,g17177);
  not NOT_6677(II25904,g17194);
  not NOT_6678(g19457,II25904);
  not NOT_6679(g19467,g16719);
  not NOT_6680(g19468,g17216);
  not NOT_6681(g19471,g18102);
  not NOT_6682(g19475,g16725);
  not NOT_6683(g19479,g16733);
  not NOT_6684(g19481,g16629);
  not NOT_6685(g19482,g17194);
  not NOT_6686(g19483,g16758);
  not NOT_6687(g19484,g16867);
  not NOT_6688(g19490,g16761);
  not NOT_6689(g19491,g17219);
  not NOT_6690(g19494,g18218);
  not NOT_6691(g19498,g16767);
  not NOT_6692(g19502,g16775);
  not NOT_6693(g19504,g16785);
  not NOT_6694(g19505,g16895);
  not NOT_6695(g19511,g16788);
  not NOT_6696(g19512,g17221);
  not NOT_6697(g19515,g18325);
  not NOT_6698(g19519,g16794);
  not NOT_6699(g19523,g16814);
  not NOT_6700(g19524,g16924);
  not NOT_6701(g19530,g16817);
  not NOT_6702(g19533,g16832);
  not NOT_6703(g19534,g16954);
  not NOT_6704(II25966,g16654);
  not NOT_6705(g19543,II25966);
  not NOT_6706(II25971,g16671);
  not NOT_6707(g19546,II25971);
  not NOT_6708(II25977,g16692);
  not NOT_6709(g19550,II25977);
  not NOT_6710(II25985,g16718);
  not NOT_6711(g19556,II25985);
  not NOT_6712(II25994,g16860);
  not NOT_6713(g19563,II25994);
  not NOT_6714(II26006,g16866);
  not NOT_6715(g19573,II26006);
  not NOT_6716(g19577,g16881);
  not NOT_6717(g19578,g16884);
  not NOT_6718(II26025,g16803);
  not NOT_6719(g19595,II26025);
  not NOT_6720(II26028,g16566);
  not NOT_6721(g19596,II26028);
  not NOT_6722(g19607,g16910);
  not NOT_6723(g19608,g16913);
  not NOT_6724(II26051,g16824);
  not NOT_6725(g19622,II26051);
  not NOT_6726(g19640,g16940);
  not NOT_6727(g19641,g16943);
  not NOT_6728(II26078,g16835);
  not NOT_6729(g19652,II26078);
  not NOT_6730(II26085,g18085);
  not NOT_6731(g19657,II26085);
  not NOT_6732(g19680,g16971);
  not NOT_6733(g19681,g16974);
  not NOT_6734(II26112,g16844);
  not NOT_6735(g19689,II26112);
  not NOT_6736(II26115,g16845);
  not NOT_6737(g19690,II26115);
  not NOT_6738(II26123,g17503);
  not NOT_6739(g19696,II26123);
  not NOT_6740(II26134,g18201);
  not NOT_6741(g19705,II26134);
  not NOT_6742(II26154,g16851);
  not NOT_6743(g19725,II26154);
  not NOT_6744(II26171,g17594);
  not NOT_6745(g19740,II26171);
  not NOT_6746(II26182,g18308);
  not NOT_6747(g19749,II26182);
  not NOT_6748(II26195,g16853);
  not NOT_6749(g19762,II26195);
  not NOT_6750(II26198,g16854);
  not NOT_6751(g19763,II26198);
  not NOT_6752(II26220,g17691);
  not NOT_6753(g19783,II26220);
  not NOT_6754(II26231,g18401);
  not NOT_6755(g19792,II26231);
  not NOT_6756(II26237,g16857);
  not NOT_6757(g19798,II26237);
  not NOT_6758(II26266,g17791);
  not NOT_6759(g19825,II26266);
  not NOT_6760(g19830,g18886);
  not NOT_6761(II26276,g16861);
  not NOT_6762(g19838,II26276);
  not NOT_6763(II26334,g18977);
  not NOT_6764(g19890,II26334);
  not NOT_6765(II26337,g16880);
  not NOT_6766(g19893,II26337);
  not NOT_6767(II26340,g17025);
  not NOT_6768(g19894,II26340);
  not NOT_6769(II26365,g18626);
  not NOT_6770(g19915,II26365);
  not NOT_6771(g19918,g18646);
  not NOT_6772(II26369,g17059);
  not NOT_6773(g19919,II26369);
  not NOT_6774(g19933,g18548);
  not NOT_6775(II26388,g17094);
  not NOT_6776(g19934,II26388);
  not NOT_6777(II26401,g17012);
  not NOT_6778(g19945,II26401);
  not NOT_6779(g19948,g17896);
  not NOT_6780(g19950,g18598);
  not NOT_6781(II26407,g17132);
  not NOT_6782(g19951,II26407);
  not NOT_6783(II26413,g16643);
  not NOT_6784(g19957,II26413);
  not NOT_6785(II26420,g17042);
  not NOT_6786(g19972,II26420);
  not NOT_6787(g19975,g18007);
  not NOT_6788(g19977,g18630);
  not NOT_6789(II26426,g16536);
  not NOT_6790(g19978,II26426);
  not NOT_6791(II26437,g16655);
  not NOT_6792(g19987,II26437);
  not NOT_6793(II26444,g17076);
  not NOT_6794(g20002,II26444);
  not NOT_6795(g20005,g18124);
  not NOT_6796(g20007,g18639);
  not NOT_6797(II26458,g17985);
  not NOT_6798(g20016,II26458);
  not NOT_6799(II26469,g16672);
  not NOT_6800(g20025,II26469);
  not NOT_6801(II26476,g17111);
  not NOT_6802(g20040,II26476);
  not NOT_6803(g20043,g18240);
  not NOT_6804(II26481,g18590);
  not NOT_6805(g20045,II26481);
  not NOT_6806(II26494,g18102);
  not NOT_6807(g20058,II26494);
  not NOT_6808(II26505,g16693);
  not NOT_6809(g20067,II26505);
  not NOT_6810(II26512,g16802);
  not NOT_6811(g20082,II26512);
  not NOT_6812(g20083,g17968);
  not NOT_6813(II26535,g18218);
  not NOT_6814(g20099,II26535);
  not NOT_6815(II26545,g16823);
  not NOT_6816(g20105,II26545);
  not NOT_6817(II26574,g18325);
  not NOT_6818(g20124,II26574);
  not NOT_6819(g20127,g18623);
  not NOT_6820(g20140,g16830);
  not NOT_6821(g20163,g17973);
  not NOT_6822(II26612,g17645);
  not NOT_6823(g20164,II26612);
  not NOT_6824(g20178,g16842);
  not NOT_6825(g20193,g18691);
  not NOT_6826(II26642,g17746);
  not NOT_6827(g20198,II26642);
  not NOT_6828(g20212,g16848);
  not NOT_6829(g20223,g18727);
  not NOT_6830(II26664,g17847);
  not NOT_6831(g20228,II26664);
  not NOT_6832(g20242,g16852);
  not NOT_6833(g20250,g18764);
  not NOT_6834(II26679,g17959);
  not NOT_6835(g20255,II26679);
  not NOT_6836(g20269,g17230);
  not NOT_6837(g20273,g18795);
  not NOT_6838(g20278,g17237);
  not NOT_6839(g20279,g17240);
  not NOT_6840(g20281,g17243);
  not NOT_6841(g20286,g17249);
  not NOT_6842(g20287,g17252);
  not NOT_6843(g20288,g17255);
  not NOT_6844(g20289,g17259);
  not NOT_6845(g20290,g17262);
  not NOT_6846(g20292,g17265);
  not NOT_6847(II26714,g17720);
  not NOT_6848(g20295,II26714);
  not NOT_6849(g20296,g17272);
  not NOT_6850(g20297,g17275);
  not NOT_6851(g20298,g17278);
  not NOT_6852(g20302,g17282);
  not NOT_6853(g20303,g17285);
  not NOT_6854(g20304,g17288);
  not NOT_6855(g20305,g17291);
  not NOT_6856(g20306,g17294);
  not NOT_6857(g20308,g17297);
  not NOT_6858(g20311,g17304);
  not NOT_6859(g20312,g17307);
  not NOT_6860(g20313,g17310);
  not NOT_6861(g20315,g17315);
  not NOT_6862(g20316,g17318);
  not NOT_6863(g20317,g17321);
  not NOT_6864(g20321,g17324);
  not NOT_6865(g20322,g17327);
  not NOT_6866(g20323,g17330);
  not NOT_6867(g20324,g17333);
  not NOT_6868(g20325,g17336);
  not NOT_6869(g20327,g17342);
  not NOT_6870(g20328,g17345);
  not NOT_6871(g20329,g17348);
  not NOT_6872(g20330,g17354);
  not NOT_6873(g20331,g17357);
  not NOT_6874(g20332,g17360);
  not NOT_6875(g20334,g17363);
  not NOT_6876(g20335,g17366);
  not NOT_6877(g20336,g17369);
  not NOT_6878(g20340,g17372);
  not NOT_6879(g20341,g17375);
  not NOT_6880(g20342,g17378);
  not NOT_6881(g20344,g17384);
  not NOT_6882(g20345,g17387);
  not NOT_6883(g20346,g17390);
  not NOT_6884(g20347,g17399);
  not NOT_6885(g20348,g17402);
  not NOT_6886(g20349,g17405);
  not NOT_6887(g20350,g17410);
  not NOT_6888(g20351,g17413);
  not NOT_6889(g20352,g17416);
  not NOT_6890(g20354,g17419);
  not NOT_6891(g20355,g17422);
  not NOT_6892(g20356,g17425);
  not NOT_6893(II26777,g17222);
  not NOT_6894(g20360,II26777);
  not NOT_6895(g20361,g17430);
  not NOT_6896(g20362,g17433);
  not NOT_6897(g20363,g17436);
  not NOT_6898(g20364,g17439);
  not NOT_6899(g20365,g17442);
  not NOT_6900(g20366,g17451);
  not NOT_6901(g20367,g17454);
  not NOT_6902(g20368,g17457);
  not NOT_6903(g20369,g17465);
  not NOT_6904(g20370,g17468);
  not NOT_6905(g20371,g17471);
  not NOT_6906(g20372,g17476);
  not NOT_6907(g20373,g17479);
  not NOT_6908(g20374,g17482);
  not NOT_6909(II26796,g17224);
  not NOT_6910(g20377,II26796);
  not NOT_6911(g20378,g17487);
  not NOT_6912(g20379,g17490);
  not NOT_6913(g20380,g17493);
  not NOT_6914(g20381,g17496);
  not NOT_6915(g20382,g17500);
  not NOT_6916(g20383,g17503);
  not NOT_6917(g20384,g17511);
  not NOT_6918(g20385,g17514);
  not NOT_6919(g20386,g17517);
  not NOT_6920(g20387,g17520);
  not NOT_6921(g20388,g17523);
  not NOT_6922(g20389,g17531);
  not NOT_6923(g20390,g17534);
  not NOT_6924(g20391,g17537);
  not NOT_6925(g20392,g17545);
  not NOT_6926(g20393,g17548);
  not NOT_6927(g20394,g17551);
  not NOT_6928(II26816,g17225);
  not NOT_6929(g20395,II26816);
  not NOT_6930(II26819,g17226);
  not NOT_6931(g20396,II26819);
  not NOT_6932(g20397,g17557);
  not NOT_6933(g20398,g17560);
  not NOT_6934(g20399,g17563);
  not NOT_6935(g20400,g17567);
  not NOT_6936(g20401,g17570);
  not NOT_6937(g20402,g17573);
  not NOT_6938(g20403,g17579);
  not NOT_6939(g20404,g17582);
  not NOT_6940(g20405,g17585);
  not NOT_6941(g20406,g17588);
  not NOT_6942(g20407,g17591);
  not NOT_6943(g20408,g17594);
  not NOT_6944(g20409,g17601);
  not NOT_6945(g20410,g17604);
  not NOT_6946(g20411,g17607);
  not NOT_6947(g20412,g17610);
  not NOT_6948(g20413,g17613);
  not NOT_6949(g20414,g17621);
  not NOT_6950(g20415,g17624);
  not NOT_6951(g20416,g17627);
  not NOT_6952(II26843,g17228);
  not NOT_6953(g20418,II26843);
  not NOT_6954(II26846,g17229);
  not NOT_6955(g20419,II26846);
  not NOT_6956(g20420,g17637);
  not NOT_6957(g20421,g17649);
  not NOT_6958(g20422,g17655);
  not NOT_6959(g20423,g17658);
  not NOT_6960(g20424,g17661);
  not NOT_6961(g20425,g17664);
  not NOT_6962(g20426,g17667);
  not NOT_6963(g20427,g17670);
  not NOT_6964(g20428,g17676);
  not NOT_6965(g20429,g17679);
  not NOT_6966(g20430,g17682);
  not NOT_6967(g20431,g17685);
  not NOT_6968(g20432,g17688);
  not NOT_6969(g20433,g17691);
  not NOT_6970(g20434,g17698);
  not NOT_6971(g20435,g17701);
  not NOT_6972(g20436,g17704);
  not NOT_6973(g20437,g17707);
  not NOT_6974(g20438,g17710);
  not NOT_6975(II26868,g17234);
  not NOT_6976(g20439,II26868);
  not NOT_6977(II26871,g17235);
  not NOT_6978(g20440,II26871);
  not NOT_6979(II26874,g17236);
  not NOT_6980(g20441,II26874);
  not NOT_6981(g20442,g17738);
  not NOT_6982(g20443,g17749);
  not NOT_6983(g20444,g17755);
  not NOT_6984(g20445,g17758);
  not NOT_6985(g20446,g17761);
  not NOT_6986(g20447,g17764);
  not NOT_6987(g20448,g17767);
  not NOT_6988(g20449,g17770);
  not NOT_6989(g20450,g17776);
  not NOT_6990(g20451,g17779);
  not NOT_6991(g20452,g17782);
  not NOT_6992(g20453,g17785);
  not NOT_6993(g20454,g17788);
  not NOT_6994(g20455,g17791);
  not NOT_6995(g20456,g17799);
  not NOT_6996(II26892,g17246);
  not NOT_6997(g20457,II26892);
  not NOT_6998(II26895,g17247);
  not NOT_6999(g20458,II26895);
  not NOT_7000(II26898,g17248);
  not NOT_7001(g20459,II26898);
  not NOT_7002(g20461,g17839);
  not NOT_7003(g20462,g17850);
  not NOT_7004(g20463,g17856);
  not NOT_7005(g20464,g17859);
  not NOT_7006(g20465,g17862);
  not NOT_7007(g20466,g17865);
  not NOT_7008(g20467,g17868);
  not NOT_7009(g20468,g17871);
  not NOT_7010(II26910,g17269);
  not NOT_7011(g20469,II26910);
  not NOT_7012(II26913,g17270);
  not NOT_7013(g20470,II26913);
  not NOT_7014(II26916,g17271);
  not NOT_7015(g20471,II26916);
  not NOT_7016(g20476,g17951);
  not NOT_7017(g20477,g17962);
  not NOT_7018(II26923,g17302);
  not NOT_7019(g20478,II26923);
  not NOT_7020(II26926,g17303);
  not NOT_7021(g20479,II26926);
  not NOT_7022(II26931,g17340);
  not NOT_7023(g20484,II26931);
  not NOT_7024(II26934,g17341);
  not NOT_7025(g20485,II26934);
  not NOT_7026(g20490,g18166);
  not NOT_7027(II26940,g17383);
  not NOT_7028(g20491,II26940);
  not NOT_7029(g20496,g18258);
  not NOT_7030(II26947,g17429);
  not NOT_7031(g20498,II26947);
  not NOT_7032(g20500,g18278);
  not NOT_7033(g20501,g18334);
  not NOT_7034(g20504,g18355);
  not NOT_7035(g20505,g18371);
  not NOT_7036(g20507,g18351);
  not NOT_7037(II26960,g16884);
  not NOT_7038(g20513,II26960);
  not NOT_7039(g20516,g18432);
  not NOT_7040(g20517,g18450);
  not NOT_7041(g20518,g18466);
  not NOT_7042(II26966,g17051);
  not NOT_7043(g20519,II26966);
  not NOT_7044(g20526,g18446);
  not NOT_7045(II26972,g16913);
  not NOT_7046(g20531,II26972);
  not NOT_7047(g20534,g18505);
  not NOT_7048(g20535,g18523);
  not NOT_7049(g20536,g18539);
  not NOT_7050(II26980,g17086);
  not NOT_7051(g20539,II26980);
  not NOT_7052(g20545,g18519);
  not NOT_7053(II26985,g16943);
  not NOT_7054(g20550,II26985);
  not NOT_7055(g20553,g18569);
  not NOT_7056(g20554,g18587);
  not NOT_7057(II26990,g19145);
  not NOT_7058(g20555,II26990);
  not NOT_7059(II26993,g19159);
  not NOT_7060(g20556,II26993);
  not NOT_7061(II26996,g19169);
  not NOT_7062(g20557,II26996);
  not NOT_7063(II26999,g19543);
  not NOT_7064(g20558,II26999);
  not NOT_7065(II27002,g19147);
  not NOT_7066(g20559,II27002);
  not NOT_7067(II27005,g19164);
  not NOT_7068(g20560,II27005);
  not NOT_7069(II27008,g19175);
  not NOT_7070(g20561,II27008);
  not NOT_7071(II27011,g19546);
  not NOT_7072(g20562,II27011);
  not NOT_7073(II27014,g19151);
  not NOT_7074(g20563,II27014);
  not NOT_7075(II27017,g19170);
  not NOT_7076(g20564,II27017);
  not NOT_7077(II27020,g19182);
  not NOT_7078(g20565,II27020);
  not NOT_7079(II27023,g19550);
  not NOT_7080(g20566,II27023);
  not NOT_7081(II27026,g19156);
  not NOT_7082(g20567,II27026);
  not NOT_7083(II27029,g19176);
  not NOT_7084(g20568,II27029);
  not NOT_7085(II27032,g19189);
  not NOT_7086(g20569,II27032);
  not NOT_7087(II27035,g19556);
  not NOT_7088(g20570,II27035);
  not NOT_7089(II27038,g20082);
  not NOT_7090(g20571,II27038);
  not NOT_7091(II27041,g19237);
  not NOT_7092(g20572,II27041);
  not NOT_7093(II27044,g19247);
  not NOT_7094(g20573,II27044);
  not NOT_7095(II27047,g19258);
  not NOT_7096(g20574,II27047);
  not NOT_7097(II27050,g19183);
  not NOT_7098(g20575,II27050);
  not NOT_7099(II27053,g19190);
  not NOT_7100(g20576,II27053);
  not NOT_7101(II27056,g19196);
  not NOT_7102(g20577,II27056);
  not NOT_7103(II27059,g19207);
  not NOT_7104(g20578,II27059);
  not NOT_7105(II27062,g19217);
  not NOT_7106(g20579,II27062);
  not NOT_7107(II27065,g19270);
  not NOT_7108(g20580,II27065);
  not NOT_7109(II27068,g19197);
  not NOT_7110(g20581,II27068);
  not NOT_7111(II27071,g19218);
  not NOT_7112(g20582,II27071);
  not NOT_7113(II27074,g19238);
  not NOT_7114(g20583,II27074);
  not NOT_7115(II27077,g19259);
  not NOT_7116(g20584,II27077);
  not NOT_7117(II27080,g19198);
  not NOT_7118(g20585,II27080);
  not NOT_7119(II27083,g19208);
  not NOT_7120(g20586,II27083);
  not NOT_7121(II27086,g19229);
  not NOT_7122(g20587,II27086);
  not NOT_7123(II27089,g20105);
  not NOT_7124(g20588,II27089);
  not NOT_7125(II27092,g19174);
  not NOT_7126(g20589,II27092);
  not NOT_7127(II27095,g19185);
  not NOT_7128(g20590,II27095);
  not NOT_7129(II27098,g19199);
  not NOT_7130(g20591,II27098);
  not NOT_7131(II27101,g19220);
  not NOT_7132(g20592,II27101);
  not NOT_7133(II27104,g19239);
  not NOT_7134(g20593,II27104);
  not NOT_7135(II27107,g19249);
  not NOT_7136(g20594,II27107);
  not NOT_7137(II27110,g19622);
  not NOT_7138(g20595,II27110);
  not NOT_7139(II27113,g19689);
  not NOT_7140(g20596,II27113);
  not NOT_7141(II27116,g19762);
  not NOT_7142(g20597,II27116);
  not NOT_7143(II27119,g19563);
  not NOT_7144(g20598,II27119);
  not NOT_7145(II27122,g19595);
  not NOT_7146(g20599,II27122);
  not NOT_7147(II27125,g19652);
  not NOT_7148(g20600,II27125);
  not NOT_7149(II27128,g19725);
  not NOT_7150(g20601,II27128);
  not NOT_7151(II27131,g19798);
  not NOT_7152(g20602,II27131);
  not NOT_7153(II27134,g19573);
  not NOT_7154(g20603,II27134);
  not NOT_7155(II27137,g19596);
  not NOT_7156(g20604,II27137);
  not NOT_7157(II27140,g19690);
  not NOT_7158(g20605,II27140);
  not NOT_7159(II27143,g19763);
  not NOT_7160(g20606,II27143);
  not NOT_7161(II27146,g19838);
  not NOT_7162(g20607,II27146);
  not NOT_7163(II27149,g19893);
  not NOT_7164(g20608,II27149);
  not NOT_7165(II27152,g20360);
  not NOT_7166(g20609,II27152);
  not NOT_7167(II27155,g20395);
  not NOT_7168(g20610,II27155);
  not NOT_7169(II27158,g20439);
  not NOT_7170(g20611,II27158);
  not NOT_7171(II27161,g20377);
  not NOT_7172(g20612,II27161);
  not NOT_7173(II27164,g20418);
  not NOT_7174(g20613,II27164);
  not NOT_7175(II27167,g20457);
  not NOT_7176(g20614,II27167);
  not NOT_7177(II27170,g20396);
  not NOT_7178(g20615,II27170);
  not NOT_7179(II27173,g20440);
  not NOT_7180(g20616,II27173);
  not NOT_7181(II27176,g20469);
  not NOT_7182(g20617,II27176);
  not NOT_7183(II27179,g20419);
  not NOT_7184(g20618,II27179);
  not NOT_7185(II27182,g20458);
  not NOT_7186(g20619,II27182);
  not NOT_7187(II27185,g20478);
  not NOT_7188(g20620,II27185);
  not NOT_7189(II27188,g20441);
  not NOT_7190(g20621,II27188);
  not NOT_7191(II27191,g20470);
  not NOT_7192(g20622,II27191);
  not NOT_7193(II27194,g20484);
  not NOT_7194(g20623,II27194);
  not NOT_7195(II27197,g20459);
  not NOT_7196(g20624,II27197);
  not NOT_7197(II27200,g20479);
  not NOT_7198(g20625,II27200);
  not NOT_7199(II27203,g20491);
  not NOT_7200(g20626,II27203);
  not NOT_7201(II27206,g20471);
  not NOT_7202(g20627,II27206);
  not NOT_7203(II27209,g20485);
  not NOT_7204(g20628,II27209);
  not NOT_7205(II27212,g20498);
  not NOT_7206(g20629,II27212);
  not NOT_7207(II27215,g19158);
  not NOT_7208(g20630,II27215);
  not NOT_7209(II27218,g19168);
  not NOT_7210(g20631,II27218);
  not NOT_7211(II27221,g19180);
  not NOT_7212(g20632,II27221);
  not NOT_7213(II27225,g19358);
  not NOT_7214(g20634,II27225);
  not NOT_7215(II27228,g19390);
  not NOT_7216(g20637,II27228);
  not NOT_7217(II27232,g19401);
  not NOT_7218(g20641,II27232);
  not NOT_7219(II27235,g19420);
  not NOT_7220(g20644,II27235);
  not NOT_7221(II27240,g19335);
  not NOT_7222(g20649,II27240);
  not NOT_7223(II27243,g19335);
  not NOT_7224(g20652,II27243);
  not NOT_7225(II27246,g19335);
  not NOT_7226(g20655,II27246);
  not NOT_7227(II27250,g19390);
  not NOT_7228(g20659,II27250);
  not NOT_7229(II27253,g19420);
  not NOT_7230(g20662,II27253);
  not NOT_7231(II27257,g19431);
  not NOT_7232(g20666,II27257);
  not NOT_7233(II27260,g19457);
  not NOT_7234(g20669,II27260);
  not NOT_7235(II27264,g19358);
  not NOT_7236(g20673,II27264);
  not NOT_7237(II27267,g19358);
  not NOT_7238(g20676,II27267);
  not NOT_7239(II27270,g19335);
  not NOT_7240(g20679,II27270);
  not NOT_7241(II27275,g19369);
  not NOT_7242(g20684,II27275);
  not NOT_7243(II27278,g19369);
  not NOT_7244(g20687,II27278);
  not NOT_7245(II27281,g19369);
  not NOT_7246(g20690,II27281);
  not NOT_7247(II27285,g19420);
  not NOT_7248(g20694,II27285);
  not NOT_7249(II27288,g19457);
  not NOT_7250(g20697,II27288);
  not NOT_7251(II27293,g19335);
  not NOT_7252(g20704,II27293);
  not NOT_7253(II27297,g19390);
  not NOT_7254(g20708,II27297);
  not NOT_7255(II27300,g19390);
  not NOT_7256(g20711,II27300);
  not NOT_7257(II27303,g19369);
  not NOT_7258(g20714,II27303);
  not NOT_7259(II27308,g19401);
  not NOT_7260(g20719,II27308);
  not NOT_7261(II27311,g19401);
  not NOT_7262(g20722,II27311);
  not NOT_7263(II27314,g19401);
  not NOT_7264(g20725,II27314);
  not NOT_7265(II27318,g19457);
  not NOT_7266(g20729,II27318);
  not NOT_7267(II27321,g19335);
  not NOT_7268(g20732,II27321);
  not NOT_7269(II27324,g19358);
  not NOT_7270(g20735,II27324);
  not NOT_7271(II27328,g19369);
  not NOT_7272(g20739,II27328);
  not NOT_7273(II27332,g19420);
  not NOT_7274(g20743,II27332);
  not NOT_7275(II27335,g19420);
  not NOT_7276(g20746,II27335);
  not NOT_7277(II27338,g19401);
  not NOT_7278(g20749,II27338);
  not NOT_7279(II27343,g19431);
  not NOT_7280(g20754,II27343);
  not NOT_7281(II27346,g19431);
  not NOT_7282(g20757,II27346);
  not NOT_7283(II27349,g19431);
  not NOT_7284(g20760,II27349);
  not NOT_7285(II27352,g19358);
  not NOT_7286(g20763,II27352);
  not NOT_7287(II27355,g19335);
  not NOT_7288(g20766,II27355);
  not NOT_7289(II27358,g19369);
  not NOT_7290(g20769,II27358);
  not NOT_7291(II27361,g19390);
  not NOT_7292(g20772,II27361);
  not NOT_7293(II27365,g19401);
  not NOT_7294(g20776,II27365);
  not NOT_7295(II27369,g19457);
  not NOT_7296(g20780,II27369);
  not NOT_7297(II27372,g19457);
  not NOT_7298(g20783,II27372);
  not NOT_7299(II27375,g19431);
  not NOT_7300(g20786,II27375);
  not NOT_7301(II27379,g19358);
  not NOT_7302(g20790,II27379);
  not NOT_7303(II27382,g19390);
  not NOT_7304(g20793,II27382);
  not NOT_7305(II27385,g19369);
  not NOT_7306(g20796,II27385);
  not NOT_7307(II27388,g19401);
  not NOT_7308(g20799,II27388);
  not NOT_7309(II27391,g19420);
  not NOT_7310(g20802,II27391);
  not NOT_7311(II27395,g19431);
  not NOT_7312(g20806,II27395);
  not NOT_7313(II27399,g19390);
  not NOT_7314(g20810,II27399);
  not NOT_7315(II27402,g19420);
  not NOT_7316(g20813,II27402);
  not NOT_7317(II27405,g19401);
  not NOT_7318(g20816,II27405);
  not NOT_7319(II27408,g19431);
  not NOT_7320(g20819,II27408);
  not NOT_7321(II27411,g19457);
  not NOT_7322(g20822,II27411);
  not NOT_7323(II27416,g19420);
  not NOT_7324(g20827,II27416);
  not NOT_7325(II27419,g19457);
  not NOT_7326(g20830,II27419);
  not NOT_7327(II27422,g19431);
  not NOT_7328(g20833,II27422);
  not NOT_7329(II27426,g19457);
  not NOT_7330(g20837,II27426);
  not NOT_7331(g20842,g19441);
  not NOT_7332(g20850,g19468);
  not NOT_7333(g20858,g19491);
  not NOT_7334(g20866,g19512);
  not NOT_7335(g20885,g19865);
  not NOT_7336(g20904,g19896);
  not NOT_7337(g20928,g19921);
  not NOT_7338(II27488,g20310);
  not NOT_7339(g20942,II27488);
  not NOT_7340(II27491,g20314);
  not NOT_7341(g20943,II27491);
  not NOT_7342(g20956,g19936);
  not NOT_7343(II27516,g20333);
  not NOT_7344(g20971,II27516);
  not NOT_7345(II27531,g20343);
  not NOT_7346(g20984,II27531);
  not NOT_7347(II27534,g20083);
  not NOT_7348(g20985,II27534);
  not NOT_7349(II27537,g19957);
  not NOT_7350(g20986,II27537);
  not NOT_7351(II27549,g20353);
  not NOT_7352(g20998,II27549);
  not NOT_7353(II27565,g19987);
  not NOT_7354(g21012,II27565);
  not NOT_7355(II27577,g20375);
  not NOT_7356(g21024,II27577);
  not NOT_7357(II27585,g20376);
  not NOT_7358(g21030,II27585);
  not NOT_7359(II27593,g20025);
  not NOT_7360(g21036,II27593);
  not NOT_7361(g21050,g20513);
  not NOT_7362(II27614,g20067);
  not NOT_7363(g21057,II27614);
  not NOT_7364(II27621,g20417);
  not NOT_7365(g21064,II27621);
  not NOT_7366(g21066,g20519);
  not NOT_7367(g21069,g20531);
  not NOT_7368(g21076,g20539);
  not NOT_7369(g21079,g20550);
  not NOT_7370(II27646,g20507);
  not NOT_7371(g21087,II27646);
  not NOT_7372(g21090,g19064);
  not NOT_7373(g21093,g19075);
  not NOT_7374(II27658,g20526);
  not NOT_7375(g21099,II27658);
  not NOT_7376(g21102,g19081);
  not NOT_7377(II27667,g20507);
  not NOT_7378(g21108,II27667);
  not NOT_7379(II27672,g20545);
  not NOT_7380(g21113,II27672);
  not NOT_7381(II27684,g20526);
  not NOT_7382(g21125,II27684);
  not NOT_7383(II27689,g19070);
  not NOT_7384(g21130,II27689);
  not NOT_7385(II27705,g20545);
  not NOT_7386(g21144,II27705);
  not NOT_7387(II27727,g19070);
  not NOT_7388(g21164,II27727);
  not NOT_7389(II27749,g19954);
  not NOT_7390(g21184,II27749);
  not NOT_7391(g21187,g19113);
  not NOT_7392(II27766,g19984);
  not NOT_7393(g21199,II27766);
  not NOT_7394(g21202,g19118);
  not NOT_7395(II27779,g20022);
  not NOT_7396(g21214,II27779);
  not NOT_7397(g21217,g19125);
  not NOT_7398(II27785,g20064);
  not NOT_7399(g21222,II27785);
  not NOT_7400(g21225,g19132);
  not NOT_7401(g21241,g19945);
  not NOT_7402(g21249,g19972);
  not NOT_7403(g21258,g20002);
  not NOT_7404(g21266,g20040);
  not NOT_7405(II27822,g19865);
  not NOT_7406(g21271,II27822);
  not NOT_7407(II27827,g19896);
  not NOT_7408(g21278,II27827);
  not NOT_7409(II27832,g19921);
  not NOT_7410(g21285,II27832);
  not NOT_7411(II27838,g19936);
  not NOT_7412(g21293,II27838);
  not NOT_7413(II27868,g19144);
  not NOT_7414(g21327,II27868);
  not NOT_7415(II27897,g19149);
  not NOT_7416(g21358,II27897);
  not NOT_7417(II27900,g19096);
  not NOT_7418(g21359,II27900);
  not NOT_7419(II27917,g19153);
  not NOT_7420(g21376,II27917);
  not NOT_7421(II27920,g19154);
  not NOT_7422(g21377,II27920);
  not NOT_7423(II27927,g19957);
  not NOT_7424(g21382,II27927);
  not NOT_7425(II27942,g19157);
  not NOT_7426(g21399,II27942);
  not NOT_7427(g21400,g19918);
  not NOT_7428(II27949,g19957);
  not NOT_7429(g21404,II27949);
  not NOT_7430(II27958,g19987);
  not NOT_7431(g21415,II27958);
  not NOT_7432(II27969,g19162);
  not NOT_7433(g21426,II27969);
  not NOT_7434(II27972,g19163);
  not NOT_7435(g21427,II27972);
  not NOT_7436(II27976,g19957);
  not NOT_7437(g21429,II27976);
  not NOT_7438(II27984,g19987);
  not NOT_7439(g21441,II27984);
  not NOT_7440(II27992,g20025);
  not NOT_7441(g21449,II27992);
  not NOT_7442(II28000,g19167);
  not NOT_7443(g21457,II28000);
  not NOT_7444(II28003,g19957);
  not NOT_7445(g21458,II28003);
  not NOT_7446(g21461,g19957);
  not NOT_7447(II28009,g20473);
  not NOT_7448(g21473,II28009);
  not NOT_7449(II28013,g19987);
  not NOT_7450(g21477,II28013);
  not NOT_7451(II28019,g20025);
  not NOT_7452(g21483,II28019);
  not NOT_7453(II28027,g20067);
  not NOT_7454(g21491,II28027);
  not NOT_7455(II28031,g19172);
  not NOT_7456(g21495,II28031);
  not NOT_7457(II28034,g19173);
  not NOT_7458(g21496,II28034);
  not NOT_7459(II28038,g19957);
  not NOT_7460(g21498,II28038);
  not NOT_7461(II28043,g19987);
  not NOT_7462(g21505,II28043);
  not NOT_7463(g21508,g19987);
  not NOT_7464(II28047,g20481);
  not NOT_7465(g21514,II28047);
  not NOT_7466(II28051,g20025);
  not NOT_7467(g21518,II28051);
  not NOT_7468(II28057,g20067);
  not NOT_7469(g21524,II28057);
  not NOT_7470(II28061,g19178);
  not NOT_7471(g21528,II28061);
  not NOT_7472(g21529,g19272);
  not NOT_7473(II28065,g19957);
  not NOT_7474(g21530,II28065);
  not NOT_7475(II28072,g19987);
  not NOT_7476(g21537,II28072);
  not NOT_7477(II28076,g20025);
  not NOT_7478(g21541,II28076);
  not NOT_7479(g21544,g20025);
  not NOT_7480(II28080,g20487);
  not NOT_7481(g21550,II28080);
  not NOT_7482(II28084,g20067);
  not NOT_7483(g21554,II28084);
  not NOT_7484(II28087,g19184);
  not NOT_7485(g21557,II28087);
  not NOT_7486(II28090,g20008);
  not NOT_7487(g21558,II28090);
  not NOT_7488(II28093,g19957);
  not NOT_7489(g21561,II28093);
  not NOT_7490(g21565,g19291);
  not NOT_7491(II28100,g19987);
  not NOT_7492(g21566,II28100);
  not NOT_7493(II28107,g20025);
  not NOT_7494(g21573,II28107);
  not NOT_7495(II28111,g20067);
  not NOT_7496(g21577,II28111);
  not NOT_7497(g21580,g20067);
  not NOT_7498(II28115,g20493);
  not NOT_7499(g21586,II28115);
  not NOT_7500(II28119,g19957);
  not NOT_7501(g21590,II28119);
  not NOT_7502(II28123,g19987);
  not NOT_7503(g21594,II28123);
  not NOT_7504(g21598,g19309);
  not NOT_7505(II28130,g20025);
  not NOT_7506(g21599,II28130);
  not NOT_7507(II28137,g20067);
  not NOT_7508(g21606,II28137);
  not NOT_7509(II28143,g19957);
  not NOT_7510(g21612,II28143);
  not NOT_7511(II28148,g19987);
  not NOT_7512(g21619,II28148);
  not NOT_7513(II28152,g20025);
  not NOT_7514(g21623,II28152);
  not NOT_7515(g21627,g19330);
  not NOT_7516(II28159,g20067);
  not NOT_7517(g21628,II28159);
  not NOT_7518(II28169,g19987);
  not NOT_7519(g21640,II28169);
  not NOT_7520(II28174,g20025);
  not NOT_7521(g21647,II28174);
  not NOT_7522(II28178,g20067);
  not NOT_7523(g21651,II28178);
  not NOT_7524(II28184,g19103);
  not NOT_7525(g21655,II28184);
  not NOT_7526(g21661,g19091);
  not NOT_7527(II28201,g20025);
  not NOT_7528(g21671,II28201);
  not NOT_7529(II28206,g20067);
  not NOT_7530(g21678,II28206);
  not NOT_7531(II28210,g20537);
  not NOT_7532(g21682,II28210);
  not NOT_7533(g21690,g19098);
  not NOT_7534(II28229,g20067);
  not NOT_7535(g21700,II28229);
  not NOT_7536(II28235,g20153);
  not NOT_7537(g21708,II28235);
  not NOT_7538(g21716,g19894);
  not NOT_7539(g21726,g19105);
  not NOT_7540(g21742,g19919);
  not NOT_7541(g21752,g19110);
  not NOT_7542(g21766,g19934);
  not NOT_7543(g21782,g19951);
  not NOT_7544(II28314,g19152);
  not NOT_7545(g21795,II28314);
  not NOT_7546(II28357,g20497);
  not NOT_7547(g21824,II28357);
  not NOT_7548(II28360,g20163);
  not NOT_7549(g21825,II28360);
  not NOT_7550(g21861,g19657);
  not NOT_7551(g21867,g19705);
  not NOT_7552(g21872,g19749);
  not NOT_7553(g21876,g19792);
  not NOT_7554(g21883,g19890);
  not NOT_7555(g21886,g19915);
  not NOT_7556(g21895,g19945);
  not NOT_7557(g21902,g19978);
  not NOT_7558(g21907,g19972);
  not NOT_7559(II28432,g19335);
  not NOT_7560(g21914,II28432);
  not NOT_7561(II28435,g19358);
  not NOT_7562(g21917,II28435);
  not NOT_7563(g21921,g20002);
  not NOT_7564(g21927,g20045);
  not NOT_7565(II28443,g19358);
  not NOT_7566(g21928,II28443);
  not NOT_7567(II28447,g19369);
  not NOT_7568(g21932,II28447);
  not NOT_7569(II28450,g19390);
  not NOT_7570(g21935,II28450);
  not NOT_7571(g21939,g20040);
  not NOT_7572(II28455,g20943);
  not NOT_7573(g21943,II28455);
  not NOT_7574(II28458,g20971);
  not NOT_7575(g21944,II28458);
  not NOT_7576(II28461,g20998);
  not NOT_7577(g21945,II28461);
  not NOT_7578(II28464,g21024);
  not NOT_7579(g21946,II28464);
  not NOT_7580(II28467,g20942);
  not NOT_7581(g21947,II28467);
  not NOT_7582(II28470,g20984);
  not NOT_7583(g21948,II28470);
  not NOT_7584(II28473,g21030);
  not NOT_7585(g21949,II28473);
  not NOT_7586(II28476,g21064);
  not NOT_7587(g21950,II28476);
  not NOT_7588(II28479,g21795);
  not NOT_7589(g21951,II28479);
  not NOT_7590(II28482,g21376);
  not NOT_7591(g21952,II28482);
  not NOT_7592(II28485,g21426);
  not NOT_7593(g21953,II28485);
  not NOT_7594(II28488,g21495);
  not NOT_7595(g21954,II28488);
  not NOT_7596(II28491,g21327);
  not NOT_7597(g21955,II28491);
  not NOT_7598(II28494,g21358);
  not NOT_7599(g21956,II28494);
  not NOT_7600(II28497,g21399);
  not NOT_7601(g21957,II28497);
  not NOT_7602(II28500,g21457);
  not NOT_7603(g21958,II28500);
  not NOT_7604(II28503,g21528);
  not NOT_7605(g21959,II28503);
  not NOT_7606(II28506,g21377);
  not NOT_7607(g21960,II28506);
  not NOT_7608(II28509,g21427);
  not NOT_7609(g21961,II28509);
  not NOT_7610(II28512,g21496);
  not NOT_7611(g21962,II28512);
  not NOT_7612(II28515,g21557);
  not NOT_7613(g21963,II28515);
  not NOT_7614(II28518,g20985);
  not NOT_7615(g21964,II28518);
  not NOT_7616(II28521,g21824);
  not NOT_7617(g21965,II28521);
  not NOT_7618(II28524,g21359);
  not NOT_7619(g21966,II28524);
  not NOT_7620(II28527,g21407);
  not NOT_7621(g21967,II28527);
  not NOT_7622(II28541,g21467);
  not NOT_7623(g21982,II28541);
  not NOT_7624(II28550,g21432);
  not NOT_7625(g21995,II28550);
  not NOT_7626(II28557,g21407);
  not NOT_7627(g22003,II28557);
  not NOT_7628(II28564,g21385);
  not NOT_7629(g22014,II28564);
  not NOT_7630(II28628,g21842);
  not NOT_7631(g22082,II28628);
  not NOT_7632(II28649,g21843);
  not NOT_7633(g22107,II28649);
  not NOT_7634(II28671,g21845);
  not NOT_7635(g22133,II28671);
  not NOT_7636(II28693,g21847);
  not NOT_7637(g22156,II28693);
  not NOT_7638(II28712,g21851);
  not NOT_7639(g22176,II28712);
  not NOT_7640(g22212,g21914);
  not NOT_7641(g22213,g21917);
  not NOT_7642(g22217,g21928);
  not NOT_7643(II28781,g21331);
  not NOT_7644(g22219,II28781);
  not NOT_7645(g22221,g21932);
  not NOT_7646(g22222,g21935);
  not NOT_7647(II28789,g21878);
  not NOT_7648(g22225,II28789);
  not NOT_7649(II28792,g21880);
  not NOT_7650(g22226,II28792);
  not NOT_7651(g22230,g20634);
  not NOT_7652(II28800,g21316);
  not NOT_7653(g22232,II28800);
  not NOT_7654(g22233,g20637);
  not NOT_7655(g22236,g20641);
  not NOT_7656(g22237,g20644);
  not NOT_7657(g22239,g20649);
  not NOT_7658(g22240,g20652);
  not NOT_7659(g22241,g20655);
  not NOT_7660(II28813,g21502);
  not NOT_7661(g22243,II28813);
  not NOT_7662(g22246,g20659);
  not NOT_7663(g22248,g20662);
  not NOT_7664(g22251,g20666);
  not NOT_7665(g22252,g20669);
  not NOT_7666(II28825,g21882);
  not NOT_7667(g22253,II28825);
  not NOT_7668(g22256,g20673);
  not NOT_7669(g22257,g20676);
  not NOT_7670(g22258,g20679);
  not NOT_7671(II28833,g21470);
  not NOT_7672(g22259,II28833);
  not NOT_7673(g22260,g20684);
  not NOT_7674(g22261,g20687);
  not NOT_7675(g22262,g20690);
  not NOT_7676(g22266,g20694);
  not NOT_7677(g22268,g20697);
  not NOT_7678(g22271,g20704);
  not NOT_7679(g22274,g20708);
  not NOT_7680(g22275,g20711);
  not NOT_7681(g22276,g20714);
  not NOT_7682(g22277,g20719);
  not NOT_7683(g22278,g20722);
  not NOT_7684(g22279,g20725);
  not NOT_7685(g22283,g20729);
  not NOT_7686(g22286,g20732);
  not NOT_7687(g22287,g20735);
  not NOT_7688(g22290,g20739);
  not NOT_7689(g22293,g20743);
  not NOT_7690(g22294,g20746);
  not NOT_7691(g22295,g20749);
  not NOT_7692(g22296,g20754);
  not NOT_7693(g22297,g20757);
  not NOT_7694(g22298,g20760);
  not NOT_7695(II28876,g21238);
  not NOT_7696(g22300,II28876);
  not NOT_7697(g22303,g20763);
  not NOT_7698(g22304,g20766);
  not NOT_7699(g22306,g20769);
  not NOT_7700(g22307,g20772);
  not NOT_7701(g22310,g20776);
  not NOT_7702(g22313,g20780);
  not NOT_7703(g22314,g20783);
  not NOT_7704(g22315,g20786);
  not NOT_7705(g22316,g21149);
  not NOT_7706(g22318,g20790);
  not NOT_7707(g22319,g21228);
  not NOT_7708(II28896,g21246);
  not NOT_7709(g22328,II28896);
  not NOT_7710(g22331,g20793);
  not NOT_7711(g22332,g20796);
  not NOT_7712(g22334,g20799);
  not NOT_7713(g22335,g20802);
  not NOT_7714(g22338,g20806);
  not NOT_7715(g22341,g21169);
  not NOT_7716(g22343,g20810);
  not NOT_7717(g22344,g21233);
  not NOT_7718(II28913,g21255);
  not NOT_7719(g22353,II28913);
  not NOT_7720(g22356,g20813);
  not NOT_7721(g22357,g20816);
  not NOT_7722(g22359,g20819);
  not NOT_7723(g22360,g20822);
  not NOT_7724(g22364,g21189);
  not NOT_7725(g22366,g20827);
  not NOT_7726(g22367,g21242);
  not NOT_7727(II28928,g21263);
  not NOT_7728(g22376,II28928);
  not NOT_7729(g22379,g20830);
  not NOT_7730(g22380,g20833);
  not NOT_7731(g22384,g21204);
  not NOT_7732(g22386,g20837);
  not NOT_7733(g22387,g21250);
  not NOT_7734(g22401,g21533);
  not NOT_7735(g22402,g21569);
  not NOT_7736(g22403,g21602);
  not NOT_7737(g22404,g21631);
  not NOT_7738(II28949,g21685);
  not NOT_7739(g22405,II28949);
  not NOT_7740(g22408,g20986);
  not NOT_7741(II28953,g21659);
  not NOT_7742(g22409,II28953);
  not NOT_7743(II28956,g21714);
  not NOT_7744(g22412,II28956);
  not NOT_7745(II28959,g21636);
  not NOT_7746(g22415,II28959);
  not NOT_7747(II28962,g21721);
  not NOT_7748(g22418,II28962);
  not NOT_7749(g22421,g21012);
  not NOT_7750(II28966,g20633);
  not NOT_7751(g22422,II28966);
  not NOT_7752(II28969,g21686);
  not NOT_7753(g22425,II28969);
  not NOT_7754(II28972,g21736);
  not NOT_7755(g22428,II28972);
  not NOT_7756(II28975,g21688);
  not NOT_7757(g22431,II28975);
  not NOT_7758(II28978,g21740);
  not NOT_7759(g22434,II28978);
  not NOT_7760(II28981,g21667);
  not NOT_7761(g22437,II28981);
  not NOT_7762(II28984,g21747);
  not NOT_7763(g22440,II28984);
  not NOT_7764(g22443,g21036);
  not NOT_7765(II28988,g20874);
  not NOT_7766(g22444,II28988);
  not NOT_7767(II28991,g20648);
  not NOT_7768(g22445,II28991);
  not NOT_7769(II28994,g21715);
  not NOT_7770(g22448,II28994);
  not NOT_7771(II28997,g21759);
  not NOT_7772(g22451,II28997);
  not NOT_7773(II29001,g20658);
  not NOT_7774(g22455,II29001);
  not NOT_7775(II29004,g21722);
  not NOT_7776(g22458,II29004);
  not NOT_7777(II29007,g21760);
  not NOT_7778(g22461,II29007);
  not NOT_7779(II29010,g21724);
  not NOT_7780(g22464,II29010);
  not NOT_7781(II29013,g21764);
  not NOT_7782(g22467,II29013);
  not NOT_7783(II29016,g21696);
  not NOT_7784(g22470,II29016);
  not NOT_7785(II29019,g21771);
  not NOT_7786(g22473,II29019);
  not NOT_7787(g22476,g21057);
  not NOT_7788(II29023,g20672);
  not NOT_7789(g22477,II29023);
  not NOT_7790(II29026,g21737);
  not NOT_7791(g22480,II29026);
  not NOT_7792(II29030,g20683);
  not NOT_7793(g22484,II29030);
  not NOT_7794(II29033,g21741);
  not NOT_7795(g22487,II29033);
  not NOT_7796(II29036,g21775);
  not NOT_7797(g22490,II29036);
  not NOT_7798(II29040,g20693);
  not NOT_7799(g22494,II29040);
  not NOT_7800(II29043,g21748);
  not NOT_7801(g22497,II29043);
  not NOT_7802(II29046,g21776);
  not NOT_7803(g22500,II29046);
  not NOT_7804(II29049,g21750);
  not NOT_7805(g22503,II29049);
  not NOT_7806(II29052,g21780);
  not NOT_7807(g22506,II29052);
  not NOT_7808(II29055,g21732);
  not NOT_7809(g22509,II29055);
  not NOT_7810(II29058,g20703);
  not NOT_7811(g22512,II29058);
  not NOT_7812(II29064,g20875);
  not NOT_7813(g22518,II29064);
  not NOT_7814(II29067,g20876);
  not NOT_7815(g22519,II29067);
  not NOT_7816(II29070,g20707);
  not NOT_7817(g22520,II29070);
  not NOT_7818(II29073,g21761);
  not NOT_7819(g22523,II29073);
  not NOT_7820(II29077,g20718);
  not NOT_7821(g22527,II29077);
  not NOT_7822(II29080,g21765);
  not NOT_7823(g22530,II29080);
  not NOT_7824(II29083,g21790);
  not NOT_7825(g22533,II29083);
  not NOT_7826(II29087,g20728);
  not NOT_7827(g22537,II29087);
  not NOT_7828(II29090,g21772);
  not NOT_7829(g22540,II29090);
  not NOT_7830(II29093,g21791);
  not NOT_7831(g22543,II29093);
  not NOT_7832(g22547,g21087);
  not NOT_7833(II29098,g20879);
  not NOT_7834(g22548,II29098);
  not NOT_7835(II29101,g20880);
  not NOT_7836(g22549,II29101);
  not NOT_7837(II29104,g20881);
  not NOT_7838(g22550,II29104);
  not NOT_7839(II29107,g21435);
  not NOT_7840(g22551,II29107);
  not NOT_7841(II29110,g20738);
  not NOT_7842(g22552,II29110);
  not NOT_7843(II29116,g20882);
  not NOT_7844(g22558,II29116);
  not NOT_7845(II29119,g20883);
  not NOT_7846(g22559,II29119);
  not NOT_7847(II29122,g20742);
  not NOT_7848(g22560,II29122);
  not NOT_7849(II29125,g21777);
  not NOT_7850(g22563,II29125);
  not NOT_7851(II29129,g20753);
  not NOT_7852(g22567,II29129);
  not NOT_7853(II29132,g21781);
  not NOT_7854(g22570,II29132);
  not NOT_7855(II29135,g21804);
  not NOT_7856(g22573,II29135);
  not NOT_7857(II29142,g20682);
  not NOT_7858(g22582,II29142);
  not NOT_7859(II29145,g20891);
  not NOT_7860(g22583,II29145);
  not NOT_7861(II29148,g20892);
  not NOT_7862(g22584,II29148);
  not NOT_7863(II29151,g20893);
  not NOT_7864(g22585,II29151);
  not NOT_7865(II29154,g20894);
  not NOT_7866(g22586,II29154);
  not NOT_7867(g22588,g21099);
  not NOT_7868(II29159,g20896);
  not NOT_7869(g22589,II29159);
  not NOT_7870(II29162,g20897);
  not NOT_7871(g22590,II29162);
  not NOT_7872(II29165,g20898);
  not NOT_7873(g22591,II29165);
  not NOT_7874(II29168,g20775);
  not NOT_7875(g22592,II29168);
  not NOT_7876(II29174,g20899);
  not NOT_7877(g22598,II29174);
  not NOT_7878(II29177,g20900);
  not NOT_7879(g22599,II29177);
  not NOT_7880(II29180,g20779);
  not NOT_7881(g22600,II29180);
  not NOT_7882(II29183,g21792);
  not NOT_7883(g22603,II29183);
  not NOT_7884(g22609,g21108);
  not NOT_7885(II29191,g20901);
  not NOT_7886(g22611,II29191);
  not NOT_7887(II29194,g20902);
  not NOT_7888(g22612,II29194);
  not NOT_7889(II29197,g20903);
  not NOT_7890(g22613,II29197);
  not NOT_7891(II29203,g20717);
  not NOT_7892(g22619,II29203);
  not NOT_7893(II29206,g20910);
  not NOT_7894(g22620,II29206);
  not NOT_7895(II29209,g20911);
  not NOT_7896(g22621,II29209);
  not NOT_7897(II29212,g20912);
  not NOT_7898(g22622,II29212);
  not NOT_7899(II29215,g20913);
  not NOT_7900(g22623,II29215);
  not NOT_7901(g22625,g21113);
  not NOT_7902(II29220,g20915);
  not NOT_7903(g22626,II29220);
  not NOT_7904(II29223,g20916);
  not NOT_7905(g22627,II29223);
  not NOT_7906(II29226,g20917);
  not NOT_7907(g22628,II29226);
  not NOT_7908(II29229,g20805);
  not NOT_7909(g22629,II29229);
  not NOT_7910(II29235,g20918);
  not NOT_7911(g22635,II29235);
  not NOT_7912(II29238,g20919);
  not NOT_7913(g22636,II29238);
  not NOT_7914(II29243,g20921);
  not NOT_7915(g22639,II29243);
  not NOT_7916(II29246,g20922);
  not NOT_7917(g22640,II29246);
  not NOT_7918(II29249,g20923);
  not NOT_7919(g22641,II29249);
  not NOT_7920(II29252,g20924);
  not NOT_7921(g22642,II29252);
  not NOT_7922(g22645,g21125);
  not NOT_7923(II29259,g20925);
  not NOT_7924(g22647,II29259);
  not NOT_7925(II29262,g20926);
  not NOT_7926(g22648,II29262);
  not NOT_7927(II29265,g20927);
  not NOT_7928(g22649,II29265);
  not NOT_7929(II29271,g20752);
  not NOT_7930(g22655,II29271);
  not NOT_7931(II29274,g20934);
  not NOT_7932(g22656,II29274);
  not NOT_7933(II29277,g20935);
  not NOT_7934(g22657,II29277);
  not NOT_7935(II29280,g20936);
  not NOT_7936(g22658,II29280);
  not NOT_7937(II29283,g20937);
  not NOT_7938(g22659,II29283);
  not NOT_7939(g22661,g21130);
  not NOT_7940(II29288,g20939);
  not NOT_7941(g22662,II29288);
  not NOT_7942(II29291,g20940);
  not NOT_7943(g22663,II29291);
  not NOT_7944(II29294,g20941);
  not NOT_7945(g22664,II29294);
  not NOT_7946(II29301,g20944);
  not NOT_7947(g22669,II29301);
  not NOT_7948(II29304,g20945);
  not NOT_7949(g22670,II29304);
  not NOT_7950(II29307,g20946);
  not NOT_7951(g22671,II29307);
  not NOT_7952(II29310,g20947);
  not NOT_7953(g22672,II29310);
  not NOT_7954(II29313,g20948);
  not NOT_7955(g22673,II29313);
  not NOT_7956(II29317,g20949);
  not NOT_7957(g22675,II29317);
  not NOT_7958(II29320,g20950);
  not NOT_7959(g22676,II29320);
  not NOT_7960(II29323,g20951);
  not NOT_7961(g22677,II29323);
  not NOT_7962(II29326,g20952);
  not NOT_7963(g22678,II29326);
  not NOT_7964(g22681,g21144);
  not NOT_7965(II29333,g20953);
  not NOT_7966(g22683,II29333);
  not NOT_7967(II29336,g20954);
  not NOT_7968(g22684,II29336);
  not NOT_7969(II29339,g20955);
  not NOT_7970(g22685,II29339);
  not NOT_7971(II29345,g20789);
  not NOT_7972(g22691,II29345);
  not NOT_7973(II29348,g20962);
  not NOT_7974(g22692,II29348);
  not NOT_7975(II29351,g20963);
  not NOT_7976(g22693,II29351);
  not NOT_7977(II29354,g20964);
  not NOT_7978(g22694,II29354);
  not NOT_7979(II29357,g20965);
  not NOT_7980(g22695,II29357);
  not NOT_7981(II29360,g21796);
  not NOT_7982(g22696,II29360);
  not NOT_7983(II29366,g20966);
  not NOT_7984(g22702,II29366);
  not NOT_7985(II29369,g20967);
  not NOT_7986(g22703,II29369);
  not NOT_7987(II29372,g20968);
  not NOT_7988(g22704,II29372);
  not NOT_7989(II29375,g20969);
  not NOT_7990(g22705,II29375);
  not NOT_7991(II29378,g20970);
  not NOT_7992(g22706,II29378);
  not NOT_7993(II29383,g20972);
  not NOT_7994(g22709,II29383);
  not NOT_7995(II29386,g20973);
  not NOT_7996(g22710,II29386);
  not NOT_7997(II29389,g20974);
  not NOT_7998(g22711,II29389);
  not NOT_7999(II29392,g20975);
  not NOT_8000(g22712,II29392);
  not NOT_8001(II29395,g20976);
  not NOT_8002(g22713,II29395);
  not NOT_8003(II29399,g20977);
  not NOT_8004(g22715,II29399);
  not NOT_8005(II29402,g20978);
  not NOT_8006(g22716,II29402);
  not NOT_8007(II29405,g20979);
  not NOT_8008(g22717,II29405);
  not NOT_8009(II29408,g20980);
  not NOT_8010(g22718,II29408);
  not NOT_8011(g22721,g21164);
  not NOT_8012(II29415,g20981);
  not NOT_8013(g22723,II29415);
  not NOT_8014(II29418,g20982);
  not NOT_8015(g22724,II29418);
  not NOT_8016(II29421,g20983);
  not NOT_8017(g22725,II29421);
  not NOT_8018(II29426,g20989);
  not NOT_8019(g22728,II29426);
  not NOT_8020(II29429,g20990);
  not NOT_8021(g22729,II29429);
  not NOT_8022(II29432,g20991);
  not NOT_8023(g22730,II29432);
  not NOT_8024(II29435,g20992);
  not NOT_8025(g22731,II29435);
  not NOT_8026(II29439,g20993);
  not NOT_8027(g22733,II29439);
  not NOT_8028(II29442,g20994);
  not NOT_8029(g22734,II29442);
  not NOT_8030(II29445,g20995);
  not NOT_8031(g22735,II29445);
  not NOT_8032(II29448,g20996);
  not NOT_8033(g22736,II29448);
  not NOT_8034(II29451,g20997);
  not NOT_8035(g22737,II29451);
  not NOT_8036(II29456,g20999);
  not NOT_8037(g22740,II29456);
  not NOT_8038(II29459,g21000);
  not NOT_8039(g22741,II29459);
  not NOT_8040(II29462,g21001);
  not NOT_8041(g22742,II29462);
  not NOT_8042(II29465,g21002);
  not NOT_8043(g22743,II29465);
  not NOT_8044(II29468,g21003);
  not NOT_8045(g22744,II29468);
  not NOT_8046(II29472,g21004);
  not NOT_8047(g22746,II29472);
  not NOT_8048(II29475,g21005);
  not NOT_8049(g22747,II29475);
  not NOT_8050(II29478,g21006);
  not NOT_8051(g22748,II29478);
  not NOT_8052(II29481,g21007);
  not NOT_8053(g22749,II29481);
  not NOT_8054(II29484,g21903);
  not NOT_8055(g22750,II29484);
  not NOT_8056(g22753,g21184);
  not NOT_8057(II29490,g21009);
  not NOT_8058(g22756,II29490);
  not NOT_8059(II29493,g21010);
  not NOT_8060(g22757,II29493);
  not NOT_8061(II29496,g21011);
  not NOT_8062(g22758,II29496);
  not NOT_8063(II29500,g21015);
  not NOT_8064(g22760,II29500);
  not NOT_8065(II29503,g21016);
  not NOT_8066(g22761,II29503);
  not NOT_8067(II29506,g21017);
  not NOT_8068(g22762,II29506);
  not NOT_8069(II29509,g21018);
  not NOT_8070(g22763,II29509);
  not NOT_8071(II29513,g21019);
  not NOT_8072(g22765,II29513);
  not NOT_8073(II29516,g21020);
  not NOT_8074(g22766,II29516);
  not NOT_8075(II29519,g21021);
  not NOT_8076(g22767,II29519);
  not NOT_8077(II29522,g21022);
  not NOT_8078(g22768,II29522);
  not NOT_8079(II29525,g21023);
  not NOT_8080(g22769,II29525);
  not NOT_8081(II29530,g21025);
  not NOT_8082(g22772,II29530);
  not NOT_8083(II29533,g21026);
  not NOT_8084(g22773,II29533);
  not NOT_8085(II29536,g21027);
  not NOT_8086(g22774,II29536);
  not NOT_8087(II29539,g21028);
  not NOT_8088(g22775,II29539);
  not NOT_8089(II29542,g21029);
  not NOT_8090(g22776,II29542);
  not NOT_8091(g22777,g21796);
  not NOT_8092(II29547,g21031);
  not NOT_8093(g22785,II29547);
  not NOT_8094(II29550,g21032);
  not NOT_8095(g22786,II29550);
  not NOT_8096(g22787,g21199);
  not NOT_8097(II29556,g21033);
  not NOT_8098(g22790,II29556);
  not NOT_8099(II29559,g21034);
  not NOT_8100(g22791,II29559);
  not NOT_8101(II29562,g21035);
  not NOT_8102(g22792,II29562);
  not NOT_8103(II29566,g21039);
  not NOT_8104(g22794,II29566);
  not NOT_8105(II29569,g21040);
  not NOT_8106(g22795,II29569);
  not NOT_8107(II29572,g21041);
  not NOT_8108(g22796,II29572);
  not NOT_8109(II29575,g21042);
  not NOT_8110(g22797,II29575);
  not NOT_8111(II29579,g21043);
  not NOT_8112(g22799,II29579);
  not NOT_8113(II29582,g21044);
  not NOT_8114(g22800,II29582);
  not NOT_8115(II29585,g21045);
  not NOT_8116(g22801,II29585);
  not NOT_8117(II29588,g21046);
  not NOT_8118(g22802,II29588);
  not NOT_8119(II29591,g21047);
  not NOT_8120(g22803,II29591);
  not NOT_8121(g22805,g21894);
  not NOT_8122(g22806,g21615);
  not NOT_8123(II29600,g21720);
  not NOT_8124(g22812,II29600);
  not NOT_8125(II29603,g21051);
  not NOT_8126(g22824,II29603);
  not NOT_8127(II29606,g21364);
  not NOT_8128(g22825,II29606);
  not NOT_8129(II29610,g21052);
  not NOT_8130(g22827,II29610);
  not NOT_8131(II29613,g21053);
  not NOT_8132(g22828,II29613);
  not NOT_8133(g22829,g21214);
  not NOT_8134(II29619,g21054);
  not NOT_8135(g22832,II29619);
  not NOT_8136(II29622,g21055);
  not NOT_8137(g22833,II29622);
  not NOT_8138(II29625,g21056);
  not NOT_8139(g22834,II29625);
  not NOT_8140(II29629,g21060);
  not NOT_8141(g22836,II29629);
  not NOT_8142(II29632,g21061);
  not NOT_8143(g22837,II29632);
  not NOT_8144(II29635,g21062);
  not NOT_8145(g22838,II29635);
  not NOT_8146(II29638,g21063);
  not NOT_8147(g22839,II29638);
  not NOT_8148(II29641,g20825);
  not NOT_8149(g22840,II29641);
  not NOT_8150(g22843,g21889);
  not NOT_8151(g22847,g21643);
  not NOT_8152(II29653,g21746);
  not NOT_8153(g22852,II29653);
  not NOT_8154(II29656,g21070);
  not NOT_8155(g22864,II29656);
  not NOT_8156(II29660,g21071);
  not NOT_8157(g22866,II29660);
  not NOT_8158(II29663,g21072);
  not NOT_8159(g22867,II29663);
  not NOT_8160(g22868,g21222);
  not NOT_8161(II29669,g21073);
  not NOT_8162(g22871,II29669);
  not NOT_8163(II29672,g21074);
  not NOT_8164(g22872,II29672);
  not NOT_8165(II29675,g21075);
  not NOT_8166(g22873,II29675);
  not NOT_8167(g22875,g21884);
  not NOT_8168(g22882,g21674);
  not NOT_8169(II29687,g21770);
  not NOT_8170(g22887,II29687);
  not NOT_8171(II29690,g21080);
  not NOT_8172(g22899,II29690);
  not NOT_8173(II29694,g21081);
  not NOT_8174(g22901,II29694);
  not NOT_8175(II29697,g21082);
  not NOT_8176(g22902,II29697);
  not NOT_8177(II29700,g20700);
  not NOT_8178(g22903,II29700);
  not NOT_8179(g22907,g21711);
  not NOT_8180(g22917,g21703);
  not NOT_8181(II29712,g21786);
  not NOT_8182(g22922,II29712);
  not NOT_8183(II29715,g21094);
  not NOT_8184(g22934,II29715);
  not NOT_8185(II29724,g21851);
  not NOT_8186(g22945,II29724);
  not NOT_8187(II29727,g20877);
  not NOT_8188(g22948,II29727);
  not NOT_8189(g22949,g21665);
  not NOT_8190(g22954,g21739);
  not NOT_8191(g22958,g21694);
  not NOT_8192(g22962,g21763);
  not NOT_8193(g22966,g21730);
  not NOT_8194(II29736,g20884);
  not NOT_8195(g22970,II29736);
  not NOT_8196(g22971,g21779);
  not NOT_8197(g22975,g21756);
  not NOT_8198(II29741,g21346);
  not NOT_8199(g22979,II29741);
  not NOT_8200(g22980,g21794);
  not NOT_8201(g22986,g21382);
  not NOT_8202(g22988,g21404);
  not NOT_8203(g22989,g21415);
  not NOT_8204(g22991,g21429);
  not NOT_8205(g22995,g21441);
  not NOT_8206(g22996,g21449);
  not NOT_8207(g22998,g21458);
  not NOT_8208(g23001,g21473);
  not NOT_8209(g23002,g21477);
  not NOT_8210(g23006,g21483);
  not NOT_8211(g23007,g21491);
  not NOT_8212(g23008,g21498);
  not NOT_8213(g23012,g21505);
  not NOT_8214(g23015,g21514);
  not NOT_8215(g23016,g21518);
  not NOT_8216(g23020,g21524);
  not NOT_8217(g23021,g21530);
  not NOT_8218(g23024,g21537);
  not NOT_8219(g23028,g21541);
  not NOT_8220(g23031,g21550);
  not NOT_8221(g23032,g21554);
  not NOT_8222(g23036,g21558);
  not NOT_8223(g23037,g21561);
  not NOT_8224(g23038,g21566);
  not NOT_8225(g23041,g21573);
  not NOT_8226(g23045,g21577);
  not NOT_8227(g23048,g21586);
  not NOT_8228(g23049,g21590);
  not NOT_8229(II29797,g21432);
  not NOT_8230(g23050,II29797);
  not NOT_8231(II29802,g21435);
  not NOT_8232(g23055,II29802);
  not NOT_8233(g23056,g21594);
  not NOT_8234(g23057,g21599);
  not NOT_8235(g23060,g21606);
  not NOT_8236(g23064,g21612);
  not NOT_8237(II29812,g21467);
  not NOT_8238(g23065,II29812);
  not NOT_8239(II29817,g21470);
  not NOT_8240(g23068,II29817);
  not NOT_8241(g23069,g21619);
  not NOT_8242(g23074,g21623);
  not NOT_8243(g23075,g21628);
  not NOT_8244(II29827,g21502);
  not NOT_8245(g23078,II29827);
  not NOT_8246(g23079,g21640);
  not NOT_8247(g23082,g21647);
  not NOT_8248(g23087,g21651);
  not NOT_8249(g23088,g21655);
  not NOT_8250(II29841,g21316);
  not NOT_8251(g23094,II29841);
  not NOT_8252(g23095,g21671);
  not NOT_8253(g23098,g21678);
  not NOT_8254(g23103,g21682);
  not NOT_8255(II29852,g21331);
  not NOT_8256(g23105,II29852);
  not NOT_8257(g23112,g21700);
  not NOT_8258(g23115,g21708);
  not NOT_8259(II29863,g21346);
  not NOT_8260(g23116,II29863);
  not NOT_8261(II29872,g21364);
  not NOT_8262(g23125,II29872);
  not NOT_8263(II29881,g21385);
  not NOT_8264(g23134,II29881);
  not NOT_8265(g23140,g21825);
  not NOT_8266(g23141,g21825);
  not NOT_8267(g23142,g21825);
  not NOT_8268(g23143,g21825);
  not NOT_8269(g23144,g21825);
  not NOT_8270(g23145,g21825);
  not NOT_8271(g23146,g21825);
  not NOT_8272(g23147,g21825);
  not NOT_8273(II29897,g23116);
  not NOT_8274(g23148,II29897);
  not NOT_8275(II29900,g23125);
  not NOT_8276(g23149,II29900);
  not NOT_8277(II29903,g23134);
  not NOT_8278(g23150,II29903);
  not NOT_8279(II29906,g21967);
  not NOT_8280(g23151,II29906);
  not NOT_8281(II29909,g23050);
  not NOT_8282(g23152,II29909);
  not NOT_8283(II29912,g23065);
  not NOT_8284(g23153,II29912);
  not NOT_8285(II29915,g23055);
  not NOT_8286(g23154,II29915);
  not NOT_8287(II29918,g23068);
  not NOT_8288(g23155,II29918);
  not NOT_8289(II29921,g23078);
  not NOT_8290(g23156,II29921);
  not NOT_8291(II29924,g23094);
  not NOT_8292(g23157,II29924);
  not NOT_8293(II29927,g23105);
  not NOT_8294(g23158,II29927);
  not NOT_8295(II29930,g22176);
  not NOT_8296(g23159,II29930);
  not NOT_8297(II29933,g22082);
  not NOT_8298(g23160,II29933);
  not NOT_8299(II29936,g22582);
  not NOT_8300(g23161,II29936);
  not NOT_8301(II29939,g22518);
  not NOT_8302(g23162,II29939);
  not NOT_8303(II29942,g22548);
  not NOT_8304(g23163,II29942);
  not NOT_8305(II29945,g22583);
  not NOT_8306(g23164,II29945);
  not NOT_8307(II29948,g22549);
  not NOT_8308(g23165,II29948);
  not NOT_8309(II29951,g22584);
  not NOT_8310(g23166,II29951);
  not NOT_8311(II29954,g22611);
  not NOT_8312(g23167,II29954);
  not NOT_8313(II29957,g22585);
  not NOT_8314(g23168,II29957);
  not NOT_8315(II29960,g22612);
  not NOT_8316(g23169,II29960);
  not NOT_8317(II29963,g22639);
  not NOT_8318(g23170,II29963);
  not NOT_8319(II29966,g22613);
  not NOT_8320(g23171,II29966);
  not NOT_8321(II29969,g22640);
  not NOT_8322(g23172,II29969);
  not NOT_8323(II29972,g22669);
  not NOT_8324(g23173,II29972);
  not NOT_8325(II29975,g22641);
  not NOT_8326(g23174,II29975);
  not NOT_8327(II29978,g22670);
  not NOT_8328(g23175,II29978);
  not NOT_8329(II29981,g22702);
  not NOT_8330(g23176,II29981);
  not NOT_8331(II29984,g22671);
  not NOT_8332(g23177,II29984);
  not NOT_8333(II29987,g22703);
  not NOT_8334(g23178,II29987);
  not NOT_8335(II29990,g22728);
  not NOT_8336(g23179,II29990);
  not NOT_8337(II29993,g22704);
  not NOT_8338(g23180,II29993);
  not NOT_8339(II29996,g22729);
  not NOT_8340(g23181,II29996);
  not NOT_8341(II29999,g22756);
  not NOT_8342(g23182,II29999);
  not NOT_8343(II30002,g22730);
  not NOT_8344(g23183,II30002);
  not NOT_8345(II30005,g22757);
  not NOT_8346(g23184,II30005);
  not NOT_8347(II30008,g22785);
  not NOT_8348(g23185,II30008);
  not NOT_8349(II30011,g22758);
  not NOT_8350(g23186,II30011);
  not NOT_8351(II30014,g22786);
  not NOT_8352(g23187,II30014);
  not NOT_8353(II30017,g22824);
  not NOT_8354(g23188,II30017);
  not NOT_8355(II30020,g22519);
  not NOT_8356(g23189,II30020);
  not NOT_8357(II30023,g22550);
  not NOT_8358(g23190,II30023);
  not NOT_8359(II30026,g22586);
  not NOT_8360(g23191,II30026);
  not NOT_8361(II30029,g22642);
  not NOT_8362(g23192,II30029);
  not NOT_8363(II30032,g22672);
  not NOT_8364(g23193,II30032);
  not NOT_8365(II30035,g22705);
  not NOT_8366(g23194,II30035);
  not NOT_8367(II30038,g22673);
  not NOT_8368(g23195,II30038);
  not NOT_8369(II30041,g22706);
  not NOT_8370(g23196,II30041);
  not NOT_8371(II30044,g22731);
  not NOT_8372(g23197,II30044);
  not NOT_8373(II30047,g22107);
  not NOT_8374(g23198,II30047);
  not NOT_8375(II30050,g22619);
  not NOT_8376(g23199,II30050);
  not NOT_8377(II30053,g22558);
  not NOT_8378(g23200,II30053);
  not NOT_8379(II30056,g22589);
  not NOT_8380(g23201,II30056);
  not NOT_8381(II30059,g22620);
  not NOT_8382(g23202,II30059);
  not NOT_8383(II30062,g22590);
  not NOT_8384(g23203,II30062);
  not NOT_8385(II30065,g22621);
  not NOT_8386(g23204,II30065);
  not NOT_8387(II30068,g22647);
  not NOT_8388(g23205,II30068);
  not NOT_8389(II30071,g22622);
  not NOT_8390(g23206,II30071);
  not NOT_8391(II30074,g22648);
  not NOT_8392(g23207,II30074);
  not NOT_8393(II30077,g22675);
  not NOT_8394(g23208,II30077);
  not NOT_8395(II30080,g22649);
  not NOT_8396(g23209,II30080);
  not NOT_8397(II30083,g22676);
  not NOT_8398(g23210,II30083);
  not NOT_8399(II30086,g22709);
  not NOT_8400(g23211,II30086);
  not NOT_8401(II30089,g22677);
  not NOT_8402(g23212,II30089);
  not NOT_8403(II30092,g22710);
  not NOT_8404(g23213,II30092);
  not NOT_8405(II30095,g22733);
  not NOT_8406(g23214,II30095);
  not NOT_8407(II30098,g22711);
  not NOT_8408(g23215,II30098);
  not NOT_8409(II30101,g22734);
  not NOT_8410(g23216,II30101);
  not NOT_8411(II30104,g22760);
  not NOT_8412(g23217,II30104);
  not NOT_8413(II30107,g22735);
  not NOT_8414(g23218,II30107);
  not NOT_8415(II30110,g22761);
  not NOT_8416(g23219,II30110);
  not NOT_8417(II30113,g22790);
  not NOT_8418(g23220,II30113);
  not NOT_8419(II30116,g22762);
  not NOT_8420(g23221,II30116);
  not NOT_8421(II30119,g22791);
  not NOT_8422(g23222,II30119);
  not NOT_8423(II30122,g22827);
  not NOT_8424(g23223,II30122);
  not NOT_8425(II30125,g22792);
  not NOT_8426(g23224,II30125);
  not NOT_8427(II30128,g22828);
  not NOT_8428(g23225,II30128);
  not NOT_8429(II30131,g22864);
  not NOT_8430(g23226,II30131);
  not NOT_8431(II30134,g22559);
  not NOT_8432(g23227,II30134);
  not NOT_8433(II30137,g22591);
  not NOT_8434(g23228,II30137);
  not NOT_8435(II30140,g22623);
  not NOT_8436(g23229,II30140);
  not NOT_8437(II30143,g22678);
  not NOT_8438(g23230,II30143);
  not NOT_8439(II30146,g22712);
  not NOT_8440(g23231,II30146);
  not NOT_8441(II30149,g22736);
  not NOT_8442(g23232,II30149);
  not NOT_8443(II30152,g22713);
  not NOT_8444(g23233,II30152);
  not NOT_8445(II30155,g22737);
  not NOT_8446(g23234,II30155);
  not NOT_8447(II30158,g22763);
  not NOT_8448(g23235,II30158);
  not NOT_8449(II30161,g22133);
  not NOT_8450(g23236,II30161);
  not NOT_8451(II30164,g22655);
  not NOT_8452(g23237,II30164);
  not NOT_8453(II30167,g22598);
  not NOT_8454(g23238,II30167);
  not NOT_8455(II30170,g22626);
  not NOT_8456(g23239,II30170);
  not NOT_8457(II30173,g22656);
  not NOT_8458(g23240,II30173);
  not NOT_8459(II30176,g22627);
  not NOT_8460(g23241,II30176);
  not NOT_8461(II30179,g22657);
  not NOT_8462(g23242,II30179);
  not NOT_8463(II30182,g22683);
  not NOT_8464(g23243,II30182);
  not NOT_8465(II30185,g22658);
  not NOT_8466(g23244,II30185);
  not NOT_8467(II30188,g22684);
  not NOT_8468(g23245,II30188);
  not NOT_8469(II30191,g22715);
  not NOT_8470(g23246,II30191);
  not NOT_8471(II30194,g22685);
  not NOT_8472(g23247,II30194);
  not NOT_8473(II30197,g22716);
  not NOT_8474(g23248,II30197);
  not NOT_8475(II30200,g22740);
  not NOT_8476(g23249,II30200);
  not NOT_8477(II30203,g22717);
  not NOT_8478(g23250,II30203);
  not NOT_8479(II30206,g22741);
  not NOT_8480(g23251,II30206);
  not NOT_8481(II30209,g22765);
  not NOT_8482(g23252,II30209);
  not NOT_8483(II30212,g22742);
  not NOT_8484(g23253,II30212);
  not NOT_8485(II30215,g22766);
  not NOT_8486(g23254,II30215);
  not NOT_8487(II30218,g22794);
  not NOT_8488(g23255,II30218);
  not NOT_8489(II30221,g22767);
  not NOT_8490(g23256,II30221);
  not NOT_8491(II30224,g22795);
  not NOT_8492(g23257,II30224);
  not NOT_8493(II30227,g22832);
  not NOT_8494(g23258,II30227);
  not NOT_8495(II30230,g22796);
  not NOT_8496(g23259,II30230);
  not NOT_8497(II30233,g22833);
  not NOT_8498(g23260,II30233);
  not NOT_8499(II30236,g22866);
  not NOT_8500(g23261,II30236);
  not NOT_8501(II30239,g22834);
  not NOT_8502(g23262,II30239);
  not NOT_8503(II30242,g22867);
  not NOT_8504(g23263,II30242);
  not NOT_8505(II30245,g22899);
  not NOT_8506(g23264,II30245);
  not NOT_8507(II30248,g22599);
  not NOT_8508(g23265,II30248);
  not NOT_8509(II30251,g22628);
  not NOT_8510(g23266,II30251);
  not NOT_8511(II30254,g22659);
  not NOT_8512(g23267,II30254);
  not NOT_8513(II30257,g22718);
  not NOT_8514(g23268,II30257);
  not NOT_8515(II30260,g22743);
  not NOT_8516(g23269,II30260);
  not NOT_8517(II30263,g22768);
  not NOT_8518(g23270,II30263);
  not NOT_8519(II30266,g22744);
  not NOT_8520(g23271,II30266);
  not NOT_8521(II30269,g22769);
  not NOT_8522(g23272,II30269);
  not NOT_8523(II30272,g22797);
  not NOT_8524(g23273,II30272);
  not NOT_8525(II30275,g22156);
  not NOT_8526(g23274,II30275);
  not NOT_8527(II30278,g22691);
  not NOT_8528(g23275,II30278);
  not NOT_8529(II30281,g22635);
  not NOT_8530(g23276,II30281);
  not NOT_8531(II30284,g22662);
  not NOT_8532(g23277,II30284);
  not NOT_8533(II30287,g22692);
  not NOT_8534(g23278,II30287);
  not NOT_8535(II30290,g22663);
  not NOT_8536(g23279,II30290);
  not NOT_8537(II30293,g22693);
  not NOT_8538(g23280,II30293);
  not NOT_8539(II30296,g22723);
  not NOT_8540(g23281,II30296);
  not NOT_8541(II30299,g22694);
  not NOT_8542(g23282,II30299);
  not NOT_8543(II30302,g22724);
  not NOT_8544(g23283,II30302);
  not NOT_8545(II30305,g22746);
  not NOT_8546(g23284,II30305);
  not NOT_8547(II30308,g22725);
  not NOT_8548(g23285,II30308);
  not NOT_8549(II30311,g22747);
  not NOT_8550(g23286,II30311);
  not NOT_8551(II30314,g22772);
  not NOT_8552(g23287,II30314);
  not NOT_8553(II30317,g22748);
  not NOT_8554(g23288,II30317);
  not NOT_8555(II30320,g22773);
  not NOT_8556(g23289,II30320);
  not NOT_8557(II30323,g22799);
  not NOT_8558(g23290,II30323);
  not NOT_8559(II30326,g22774);
  not NOT_8560(g23291,II30326);
  not NOT_8561(II30329,g22800);
  not NOT_8562(g23292,II30329);
  not NOT_8563(II30332,g22836);
  not NOT_8564(g23293,II30332);
  not NOT_8565(II30335,g22801);
  not NOT_8566(g23294,II30335);
  not NOT_8567(II30338,g22837);
  not NOT_8568(g23295,II30338);
  not NOT_8569(II30341,g22871);
  not NOT_8570(g23296,II30341);
  not NOT_8571(II30344,g22838);
  not NOT_8572(g23297,II30344);
  not NOT_8573(II30347,g22872);
  not NOT_8574(g23298,II30347);
  not NOT_8575(II30350,g22901);
  not NOT_8576(g23299,II30350);
  not NOT_8577(II30353,g22873);
  not NOT_8578(g23300,II30353);
  not NOT_8579(II30356,g22902);
  not NOT_8580(g23301,II30356);
  not NOT_8581(II30359,g22934);
  not NOT_8582(g23302,II30359);
  not NOT_8583(II30362,g22636);
  not NOT_8584(g23303,II30362);
  not NOT_8585(II30365,g22664);
  not NOT_8586(g23304,II30365);
  not NOT_8587(II30368,g22695);
  not NOT_8588(g23305,II30368);
  not NOT_8589(II30371,g22749);
  not NOT_8590(g23306,II30371);
  not NOT_8591(II30374,g22775);
  not NOT_8592(g23307,II30374);
  not NOT_8593(II30377,g22802);
  not NOT_8594(g23308,II30377);
  not NOT_8595(II30380,g22776);
  not NOT_8596(g23309,II30380);
  not NOT_8597(II30383,g22803);
  not NOT_8598(g23310,II30383);
  not NOT_8599(II30386,g22839);
  not NOT_8600(g23311,II30386);
  not NOT_8601(II30389,g22225);
  not NOT_8602(g23312,II30389);
  not NOT_8603(II30392,g22226);
  not NOT_8604(g23313,II30392);
  not NOT_8605(II30395,g22253);
  not NOT_8606(g23314,II30395);
  not NOT_8607(II30398,g22840);
  not NOT_8608(g23315,II30398);
  not NOT_8609(II30401,g22444);
  not NOT_8610(g23316,II30401);
  not NOT_8611(II30404,g22948);
  not NOT_8612(g23317,II30404);
  not NOT_8613(II30407,g22970);
  not NOT_8614(g23318,II30407);
  not NOT_8615(g23403,g23052);
  not NOT_8616(g23410,g23071);
  not NOT_8617(g23415,g23084);
  not NOT_8618(g23420,g23089);
  not NOT_8619(g23424,g23100);
  not NOT_8620(g23429,g23107);
  not NOT_8621(g23435,g23120);
  not NOT_8622(II30467,g23000);
  not NOT_8623(g23438,II30467);
  not NOT_8624(II30470,g23117);
  not NOT_8625(g23439,II30470);
  not NOT_8626(g23441,g23129);
  not NOT_8627(g23444,g22945);
  not NOT_8628(II30476,g22876);
  not NOT_8629(g23448,II30476);
  not NOT_8630(II30480,g23014);
  not NOT_8631(g23452,II30480);
  not NOT_8632(II30483,g23126);
  not NOT_8633(g23453,II30483);
  not NOT_8634(II30486,g23022);
  not NOT_8635(g23454,II30486);
  not NOT_8636(II30489,g22911);
  not NOT_8637(g23455,II30489);
  not NOT_8638(II30493,g23030);
  not NOT_8639(g23459,II30493);
  not NOT_8640(II30496,g23137);
  not NOT_8641(g23460,II30496);
  not NOT_8642(II30501,g23039);
  not NOT_8643(g23463,II30501);
  not NOT_8644(II30504,g22936);
  not NOT_8645(g23464,II30504);
  not NOT_8646(II30508,g23047);
  not NOT_8647(g23468,II30508);
  not NOT_8648(II30511,g21970);
  not NOT_8649(g23469,II30511);
  not NOT_8650(g23470,g22188);
  not NOT_8651(II30516,g23058);
  not NOT_8652(g23472,II30516);
  not NOT_8653(II30519,g22942);
  not NOT_8654(g23473,II30519);
  not NOT_8655(II30525,g23067);
  not NOT_8656(g23481,II30525);
  not NOT_8657(g23482,g22197);
  not NOT_8658(II30531,g23076);
  not NOT_8659(g23485,II30531);
  not NOT_8660(II30536,g23081);
  not NOT_8661(g23492,II30536);
  not NOT_8662(g23493,g22203);
  not NOT_8663(II30544,g23092);
  not NOT_8664(g23500,II30544);
  not NOT_8665(II30547,g23093);
  not NOT_8666(g23501,II30547);
  not NOT_8667(II30552,g23097);
  not NOT_8668(g23508,II30552);
  not NOT_8669(g23509,g22209);
  not NOT_8670(II30560,g23110);
  not NOT_8671(g23516,II30560);
  not NOT_8672(II30563,g23111);
  not NOT_8673(g23517,II30563);
  not NOT_8674(II30568,g23114);
  not NOT_8675(g23524,II30568);
  not NOT_8676(II30575,g23123);
  not NOT_8677(g23531,II30575);
  not NOT_8678(II30578,g23124);
  not NOT_8679(g23532,II30578);
  not NOT_8680(II30586,g23132);
  not NOT_8681(g23542,II30586);
  not NOT_8682(II30589,g23133);
  not NOT_8683(g23543,II30589);
  not NOT_8684(II30594,g22025);
  not NOT_8685(g23546,II30594);
  not NOT_8686(II30598,g22027);
  not NOT_8687(g23548,II30598);
  not NOT_8688(II30601,g22028);
  not NOT_8689(g23549,II30601);
  not NOT_8690(II30607,g22029);
  not NOT_8691(g23553,II30607);
  not NOT_8692(II30611,g22030);
  not NOT_8693(g23555,II30611);
  not NOT_8694(II30614,g22031);
  not NOT_8695(g23556,II30614);
  not NOT_8696(II30617,g22032);
  not NOT_8697(g23557,II30617);
  not NOT_8698(II30623,g22033);
  not NOT_8699(g23561,II30623);
  not NOT_8700(II30626,g22034);
  not NOT_8701(g23562,II30626);
  not NOT_8702(II30632,g22035);
  not NOT_8703(g23566,II30632);
  not NOT_8704(II30636,g22037);
  not NOT_8705(g23568,II30636);
  not NOT_8706(II30639,g22038);
  not NOT_8707(g23569,II30639);
  not NOT_8708(II30642,g22039);
  not NOT_8709(g23570,II30642);
  not NOT_8710(II30648,g22040);
  not NOT_8711(g23574,II30648);
  not NOT_8712(II30651,g22041);
  not NOT_8713(g23575,II30651);
  not NOT_8714(II30654,g22042);
  not NOT_8715(g23576,II30654);
  not NOT_8716(II30660,g22043);
  not NOT_8717(g23580,II30660);
  not NOT_8718(II30663,g22044);
  not NOT_8719(g23581,II30663);
  not NOT_8720(II30669,g22045);
  not NOT_8721(g23585,II30669);
  not NOT_8722(II30673,g22047);
  not NOT_8723(g23587,II30673);
  not NOT_8724(II30676,g22048);
  not NOT_8725(g23588,II30676);
  not NOT_8726(II30679,g22049);
  not NOT_8727(g23589,II30679);
  not NOT_8728(II30686,g23136);
  not NOT_8729(g23594,II30686);
  not NOT_8730(II30689,g22054);
  not NOT_8731(g23595,II30689);
  not NOT_8732(II30692,g22055);
  not NOT_8733(g23596,II30692);
  not NOT_8734(II30695,g22056);
  not NOT_8735(g23597,II30695);
  not NOT_8736(II30701,g22057);
  not NOT_8737(g23601,II30701);
  not NOT_8738(II30704,g22058);
  not NOT_8739(g23602,II30704);
  not NOT_8740(II30707,g22059);
  not NOT_8741(g23603,II30707);
  not NOT_8742(II30713,g22060);
  not NOT_8743(g23607,II30713);
  not NOT_8744(II30716,g22061);
  not NOT_8745(g23608,II30716);
  not NOT_8746(II30722,g22063);
  not NOT_8747(g23612,II30722);
  not NOT_8748(II30725,g22064);
  not NOT_8749(g23613,II30725);
  not NOT_8750(II30728,g22065);
  not NOT_8751(g23614,II30728);
  not NOT_8752(II30735,g22066);
  not NOT_8753(g23619,II30735);
  not NOT_8754(II30738,g22067);
  not NOT_8755(g23620,II30738);
  not NOT_8756(II30741,g22068);
  not NOT_8757(g23621,II30741);
  not NOT_8758(II30748,g21969);
  not NOT_8759(g23626,II30748);
  not NOT_8760(II30751,g22073);
  not NOT_8761(g23627,II30751);
  not NOT_8762(II30754,g22074);
  not NOT_8763(g23628,II30754);
  not NOT_8764(II30757,g22075);
  not NOT_8765(g23629,II30757);
  not NOT_8766(II30763,g22076);
  not NOT_8767(g23633,II30763);
  not NOT_8768(II30766,g22077);
  not NOT_8769(g23634,II30766);
  not NOT_8770(II30769,g22078);
  not NOT_8771(g23635,II30769);
  not NOT_8772(II30776,g22079);
  not NOT_8773(g23640,II30776);
  not NOT_8774(II30779,g22080);
  not NOT_8775(g23641,II30779);
  not NOT_8776(II30782,g22081);
  not NOT_8777(g23642,II30782);
  not NOT_8778(II30786,g22454);
  not NOT_8779(g23644,II30786);
  not NOT_8780(II30797,g22087);
  not NOT_8781(g23661,II30797);
  not NOT_8782(II30800,g22088);
  not NOT_8783(g23662,II30800);
  not NOT_8784(II30803,g22089);
  not NOT_8785(g23663,II30803);
  not NOT_8786(II30810,g22090);
  not NOT_8787(g23668,II30810);
  not NOT_8788(II30813,g22091);
  not NOT_8789(g23669,II30813);
  not NOT_8790(II30816,g22092);
  not NOT_8791(g23670,II30816);
  not NOT_8792(II30823,g21972);
  not NOT_8793(g23675,II30823);
  not NOT_8794(II30826,g22097);
  not NOT_8795(g23676,II30826);
  not NOT_8796(II30829,g22098);
  not NOT_8797(g23677,II30829);
  not NOT_8798(II30832,g22099);
  not NOT_8799(g23678,II30832);
  not NOT_8800(II30838,g22100);
  not NOT_8801(g23682,II30838);
  not NOT_8802(II30841,g22101);
  not NOT_8803(g23683,II30841);
  not NOT_8804(II30844,g22102);
  not NOT_8805(g23684,II30844);
  not NOT_8806(II30847,g22103);
  not NOT_8807(g23685,II30847);
  not NOT_8808(II30854,g22104);
  not NOT_8809(g23690,II30854);
  not NOT_8810(II30857,g22105);
  not NOT_8811(g23691,II30857);
  not NOT_8812(II30860,g22106);
  not NOT_8813(g23692,II30860);
  not NOT_8814(II30864,g22493);
  not NOT_8815(g23694,II30864);
  not NOT_8816(II30875,g22112);
  not NOT_8817(g23711,II30875);
  not NOT_8818(II30878,g22113);
  not NOT_8819(g23712,II30878);
  not NOT_8820(II30881,g22114);
  not NOT_8821(g23713,II30881);
  not NOT_8822(II30888,g22115);
  not NOT_8823(g23718,II30888);
  not NOT_8824(II30891,g22116);
  not NOT_8825(g23719,II30891);
  not NOT_8826(II30894,g22117);
  not NOT_8827(g23720,II30894);
  not NOT_8828(II30901,g21974);
  not NOT_8829(g23725,II30901);
  not NOT_8830(II30905,g22122);
  not NOT_8831(g23727,II30905);
  not NOT_8832(II30908,g22123);
  not NOT_8833(g23728,II30908);
  not NOT_8834(II30911,g22124);
  not NOT_8835(g23729,II30911);
  not NOT_8836(II30914,g22125);
  not NOT_8837(g23730,II30914);
  not NOT_8838(II30917,g22806);
  not NOT_8839(g23731,II30917);
  not NOT_8840(II30922,g22126);
  not NOT_8841(g23736,II30922);
  not NOT_8842(II30925,g22127);
  not NOT_8843(g23737,II30925);
  not NOT_8844(II30928,g22128);
  not NOT_8845(g23738,II30928);
  not NOT_8846(II30931,g22129);
  not NOT_8847(g23739,II30931);
  not NOT_8848(II30938,g22130);
  not NOT_8849(g23744,II30938);
  not NOT_8850(II30941,g22131);
  not NOT_8851(g23745,II30941);
  not NOT_8852(II30944,g22132);
  not NOT_8853(g23746,II30944);
  not NOT_8854(II30948,g22536);
  not NOT_8855(g23748,II30948);
  not NOT_8856(II30959,g22138);
  not NOT_8857(g23765,II30959);
  not NOT_8858(II30962,g22139);
  not NOT_8859(g23766,II30962);
  not NOT_8860(II30965,g22140);
  not NOT_8861(g23767,II30965);
  not NOT_8862(II30973,g22141);
  not NOT_8863(g23773,II30973);
  not NOT_8864(II30976,g22142);
  not NOT_8865(g23774,II30976);
  not NOT_8866(II30979,g22143);
  not NOT_8867(g23775,II30979);
  not NOT_8868(II30985,g22992);
  not NOT_8869(g23779,II30985);
  not NOT_8870(II30988,g22145);
  not NOT_8871(g23782,II30988);
  not NOT_8872(II30991,g22146);
  not NOT_8873(g23783,II30991);
  not NOT_8874(II30994,g22147);
  not NOT_8875(g23784,II30994);
  not NOT_8876(II30997,g22148);
  not NOT_8877(g23785,II30997);
  not NOT_8878(II31000,g22847);
  not NOT_8879(g23786,II31000);
  not NOT_8880(II31005,g22149);
  not NOT_8881(g23791,II31005);
  not NOT_8882(II31008,g22150);
  not NOT_8883(g23792,II31008);
  not NOT_8884(II31011,g22151);
  not NOT_8885(g23793,II31011);
  not NOT_8886(II31014,g22152);
  not NOT_8887(g23794,II31014);
  not NOT_8888(II31021,g22153);
  not NOT_8889(g23799,II31021);
  not NOT_8890(II31024,g22154);
  not NOT_8891(g23800,II31024);
  not NOT_8892(II31027,g22155);
  not NOT_8893(g23801,II31027);
  not NOT_8894(II31031,g22576);
  not NOT_8895(g23803,II31031);
  not NOT_8896(II31043,g22161);
  not NOT_8897(g23821,II31043);
  not NOT_8898(II31050,g22162);
  not NOT_8899(g23826,II31050);
  not NOT_8900(II31053,g22163);
  not NOT_8901(g23827,II31053);
  not NOT_8902(II31056,g22164);
  not NOT_8903(g23828,II31056);
  not NOT_8904(II31062,g23003);
  not NOT_8905(g23832,II31062);
  not NOT_8906(II31065,g22166);
  not NOT_8907(g23835,II31065);
  not NOT_8908(II31068,g22167);
  not NOT_8909(g23836,II31068);
  not NOT_8910(II31071,g22168);
  not NOT_8911(g23837,II31071);
  not NOT_8912(II31074,g22169);
  not NOT_8913(g23838,II31074);
  not NOT_8914(II31077,g22882);
  not NOT_8915(g23839,II31077);
  not NOT_8916(II31082,g22170);
  not NOT_8917(g23844,II31082);
  not NOT_8918(II31085,g22171);
  not NOT_8919(g23845,II31085);
  not NOT_8920(II31088,g22172);
  not NOT_8921(g23846,II31088);
  not NOT_8922(II31091,g22173);
  not NOT_8923(g23847,II31091);
  not NOT_8924(g23853,g22300);
  not NOT_8925(II31102,g22177);
  not NOT_8926(g23856,II31102);
  not NOT_8927(II31109,g22178);
  not NOT_8928(g23861,II31109);
  not NOT_8929(II31112,g22179);
  not NOT_8930(g23862,II31112);
  not NOT_8931(II31115,g22180);
  not NOT_8932(g23863,II31115);
  not NOT_8933(II31121,g23017);
  not NOT_8934(g23867,II31121);
  not NOT_8935(II31124,g22182);
  not NOT_8936(g23870,II31124);
  not NOT_8937(II31127,g22183);
  not NOT_8938(g23871,II31127);
  not NOT_8939(II31130,g22184);
  not NOT_8940(g23872,II31130);
  not NOT_8941(II31133,g22185);
  not NOT_8942(g23873,II31133);
  not NOT_8943(II31136,g22917);
  not NOT_8944(g23874,II31136);
  not NOT_8945(II31141,g22777);
  not NOT_8946(g23879,II31141);
  not NOT_8947(II31144,g22935);
  not NOT_8948(g23882,II31144);
  not NOT_8949(g23885,g22062);
  not NOT_8950(g23887,g22328);
  not NOT_8951(II31152,g22191);
  not NOT_8952(g23890,II31152);
  not NOT_8953(II31159,g22192);
  not NOT_8954(g23895,II31159);
  not NOT_8955(II31162,g22193);
  not NOT_8956(g23896,II31162);
  not NOT_8957(II31165,g22194);
  not NOT_8958(g23897,II31165);
  not NOT_8959(II31171,g23033);
  not NOT_8960(g23901,II31171);
  not NOT_8961(g23905,g22046);
  not NOT_8962(g23908,g22353);
  not NOT_8963(II31181,g22200);
  not NOT_8964(g23911,II31181);
  not NOT_8965(II31188,g21989);
  not NOT_8966(g23916,II31188);
  not NOT_8967(g23918,g22036);
  not NOT_8968(II31195,g22578);
  not NOT_8969(g23923,II31195);
  not NOT_8970(g23940,g22376);
  not NOT_8971(II31205,g22002);
  not NOT_8972(g23943,II31205);
  not NOT_8973(II31213,g22615);
  not NOT_8974(g23955,II31213);
  not NOT_8975(II31226,g22651);
  not NOT_8976(g23984,II31226);
  not NOT_8977(II31232,g22026);
  not NOT_8978(g24000,II31232);
  not NOT_8979(II31235,g22218);
  not NOT_8980(g24001,II31235);
  not NOT_8981(II31244,g22687);
  not NOT_8982(g24014,II31244);
  not NOT_8983(II31250,g22953);
  not NOT_8984(g24030,II31250);
  not NOT_8985(II31253,g22231);
  not NOT_8986(g24033,II31253);
  not NOT_8987(II31257,g22234);
  not NOT_8988(g24035,II31257);
  not NOT_8989(g24047,g23023);
  not NOT_8990(II31266,g22242);
  not NOT_8991(g24051,II31266);
  not NOT_8992(II31270,g22247);
  not NOT_8993(g24053,II31270);
  not NOT_8994(II31274,g22249);
  not NOT_8995(g24055,II31274);
  not NOT_8996(g24060,g23040);
  not NOT_8997(II31282,g22263);
  not NOT_8998(g24064,II31282);
  not NOT_8999(II31286,g22267);
  not NOT_9000(g24066,II31286);
  not NOT_9001(II31290,g22269);
  not NOT_9002(g24068,II31290);
  not NOT_9003(g24073,g23059);
  not NOT_9004(II31298,g22280);
  not NOT_9005(g24077,II31298);
  not NOT_9006(II31302,g22284);
  not NOT_9007(g24079,II31302);
  not NOT_9008(g24084,g23077);
  not NOT_9009(II31310,g22299);
  not NOT_9010(g24088,II31310);
  not NOT_9011(g24094,g22339);
  not NOT_9012(g24095,g22362);
  not NOT_9013(g24096,g22405);
  not NOT_9014(g24097,g22382);
  not NOT_9015(g24098,g22409);
  not NOT_9016(g24099,g22412);
  not NOT_9017(g24101,g22415);
  not NOT_9018(g24102,g22418);
  not NOT_9019(g24103,g22397);
  not NOT_9020(g24104,g22422);
  not NOT_9021(g24105,g22425);
  not NOT_9022(g24106,g22428);
  not NOT_9023(g24107,g22431);
  not NOT_9024(g24108,g22434);
  not NOT_9025(g24110,g22437);
  not NOT_9026(g24111,g22440);
  not NOT_9027(g24112,g22445);
  not NOT_9028(g24113,g22448);
  not NOT_9029(g24114,g22451);
  not NOT_9030(g24115,g22381);
  not NOT_9031(g24121,g22455);
  not NOT_9032(g24122,g22458);
  not NOT_9033(g24123,g22461);
  not NOT_9034(g24124,g22464);
  not NOT_9035(g24125,g22467);
  not NOT_9036(g24127,g22470);
  not NOT_9037(g24128,g22473);
  not NOT_9038(g24129,g22477);
  not NOT_9039(g24130,g22480);
  not NOT_9040(g24131,g22484);
  not NOT_9041(g24132,g22487);
  not NOT_9042(g24133,g22490);
  not NOT_9043(g24134,g22396);
  not NOT_9044(g24140,g22494);
  not NOT_9045(g24141,g22497);
  not NOT_9046(g24142,g22500);
  not NOT_9047(g24143,g22503);
  not NOT_9048(g24144,g22506);
  not NOT_9049(g24146,g22509);
  not NOT_9050(g24147,g22512);
  not NOT_9051(g24148,g22520);
  not NOT_9052(g24149,g22523);
  not NOT_9053(g24150,g22527);
  not NOT_9054(g24151,g22530);
  not NOT_9055(g24152,g22533);
  not NOT_9056(g24153,g22399);
  not NOT_9057(g24159,g22537);
  not NOT_9058(g24160,g22540);
  not NOT_9059(g24161,g22543);
  not NOT_9060(g24162,g22552);
  not NOT_9061(g24163,g22560);
  not NOT_9062(g24164,g22563);
  not NOT_9063(g24165,g22567);
  not NOT_9064(g24166,g22570);
  not NOT_9065(g24167,g22573);
  not NOT_9066(g24168,g22400);
  not NOT_9067(g24175,g22592);
  not NOT_9068(g24176,g22600);
  not NOT_9069(g24177,g22603);
  not NOT_9070(g24180,g22629);
  not NOT_9071(II31387,g22811);
  not NOT_9072(g24183,II31387);
  not NOT_9073(g24210,g22696);
  not NOT_9074(g24220,g22750);
  not NOT_9075(II31417,g22578);
  not NOT_9076(g24233,II31417);
  not NOT_9077(II31426,g22615);
  not NOT_9078(g24240,II31426);
  not NOT_9079(II31436,g22651);
  not NOT_9080(g24248,II31436);
  not NOT_9081(g24251,g22903);
  not NOT_9082(II31445,g22687);
  not NOT_9083(g24255,II31445);
  not NOT_9084(II31451,g23682);
  not NOT_9085(g24259,II31451);
  not NOT_9086(II31454,g23727);
  not NOT_9087(g24260,II31454);
  not NOT_9088(II31457,g23773);
  not NOT_9089(g24261,II31457);
  not NOT_9090(II31460,g23728);
  not NOT_9091(g24262,II31460);
  not NOT_9092(II31463,g23774);
  not NOT_9093(g24263,II31463);
  not NOT_9094(II31466,g23821);
  not NOT_9095(g24264,II31466);
  not NOT_9096(II31469,g23546);
  not NOT_9097(g24265,II31469);
  not NOT_9098(II31472,g23548);
  not NOT_9099(g24266,II31472);
  not NOT_9100(II31475,g23555);
  not NOT_9101(g24267,II31475);
  not NOT_9102(II31478,g23549);
  not NOT_9103(g24268,II31478);
  not NOT_9104(II31481,g23556);
  not NOT_9105(g24269,II31481);
  not NOT_9106(II31484,g23568);
  not NOT_9107(g24270,II31484);
  not NOT_9108(II31487,g23557);
  not NOT_9109(g24271,II31487);
  not NOT_9110(II31490,g23569);
  not NOT_9111(g24272,II31490);
  not NOT_9112(II31493,g23587);
  not NOT_9113(g24273,II31493);
  not NOT_9114(II31496,g23570);
  not NOT_9115(g24274,II31496);
  not NOT_9116(II31499,g23588);
  not NOT_9117(g24275,II31499);
  not NOT_9118(II31502,g23612);
  not NOT_9119(g24276,II31502);
  not NOT_9120(II31505,g23589);
  not NOT_9121(g24277,II31505);
  not NOT_9122(II31508,g23613);
  not NOT_9123(g24278,II31508);
  not NOT_9124(II31511,g23640);
  not NOT_9125(g24279,II31511);
  not NOT_9126(II31514,g23614);
  not NOT_9127(g24280,II31514);
  not NOT_9128(II31517,g23641);
  not NOT_9129(g24281,II31517);
  not NOT_9130(II31520,g23683);
  not NOT_9131(g24282,II31520);
  not NOT_9132(II31523,g23642);
  not NOT_9133(g24283,II31523);
  not NOT_9134(II31526,g23684);
  not NOT_9135(g24284,II31526);
  not NOT_9136(II31529,g23729);
  not NOT_9137(g24285,II31529);
  not NOT_9138(II31532,g23685);
  not NOT_9139(g24286,II31532);
  not NOT_9140(II31535,g23730);
  not NOT_9141(g24287,II31535);
  not NOT_9142(II31538,g23775);
  not NOT_9143(g24288,II31538);
  not NOT_9144(II31541,g23500);
  not NOT_9145(g24289,II31541);
  not NOT_9146(II31544,g23438);
  not NOT_9147(g24290,II31544);
  not NOT_9148(II31547,g23454);
  not NOT_9149(g24291,II31547);
  not NOT_9150(II31550,g23481);
  not NOT_9151(g24292,II31550);
  not NOT_9152(II31553,g23501);
  not NOT_9153(g24293,II31553);
  not NOT_9154(II31556,g23439);
  not NOT_9155(g24294,II31556);
  not NOT_9156(II31559,g24233);
  not NOT_9157(g24295,II31559);
  not NOT_9158(II31562,g23594);
  not NOT_9159(g24296,II31562);
  not NOT_9160(II31565,g24001);
  not NOT_9161(g24297,II31565);
  not NOT_9162(II31568,g24033);
  not NOT_9163(g24298,II31568);
  not NOT_9164(II31571,g24051);
  not NOT_9165(g24299,II31571);
  not NOT_9166(II31574,g23736);
  not NOT_9167(g24300,II31574);
  not NOT_9168(II31577,g23782);
  not NOT_9169(g24301,II31577);
  not NOT_9170(II31580,g23826);
  not NOT_9171(g24302,II31580);
  not NOT_9172(II31583,g23783);
  not NOT_9173(g24303,II31583);
  not NOT_9174(II31586,g23827);
  not NOT_9175(g24304,II31586);
  not NOT_9176(II31589,g23856);
  not NOT_9177(g24305,II31589);
  not NOT_9178(II31592,g23553);
  not NOT_9179(g24306,II31592);
  not NOT_9180(II31595,g23561);
  not NOT_9181(g24307,II31595);
  not NOT_9182(II31598,g23574);
  not NOT_9183(g24308,II31598);
  not NOT_9184(II31601,g23562);
  not NOT_9185(g24309,II31601);
  not NOT_9186(II31604,g23575);
  not NOT_9187(g24310,II31604);
  not NOT_9188(II31607,g23595);
  not NOT_9189(g24311,II31607);
  not NOT_9190(II31610,g23576);
  not NOT_9191(g24312,II31610);
  not NOT_9192(II31613,g23596);
  not NOT_9193(g24313,II31613);
  not NOT_9194(II31616,g23619);
  not NOT_9195(g24314,II31616);
  not NOT_9196(II31619,g23597);
  not NOT_9197(g24315,II31619);
  not NOT_9198(II31622,g23620);
  not NOT_9199(g24316,II31622);
  not NOT_9200(II31625,g23661);
  not NOT_9201(g24317,II31625);
  not NOT_9202(II31628,g23621);
  not NOT_9203(g24318,II31628);
  not NOT_9204(II31631,g23662);
  not NOT_9205(g24319,II31631);
  not NOT_9206(II31634,g23690);
  not NOT_9207(g24320,II31634);
  not NOT_9208(II31637,g23663);
  not NOT_9209(g24321,II31637);
  not NOT_9210(II31640,g23691);
  not NOT_9211(g24322,II31640);
  not NOT_9212(II31643,g23737);
  not NOT_9213(g24323,II31643);
  not NOT_9214(II31646,g23692);
  not NOT_9215(g24324,II31646);
  not NOT_9216(II31649,g23738);
  not NOT_9217(g24325,II31649);
  not NOT_9218(II31652,g23784);
  not NOT_9219(g24326,II31652);
  not NOT_9220(II31655,g23739);
  not NOT_9221(g24327,II31655);
  not NOT_9222(II31658,g23785);
  not NOT_9223(g24328,II31658);
  not NOT_9224(II31661,g23828);
  not NOT_9225(g24329,II31661);
  not NOT_9226(II31664,g23516);
  not NOT_9227(g24330,II31664);
  not NOT_9228(II31667,g23452);
  not NOT_9229(g24331,II31667);
  not NOT_9230(II31670,g23463);
  not NOT_9231(g24332,II31670);
  not NOT_9232(II31673,g23492);
  not NOT_9233(g24333,II31673);
  not NOT_9234(II31676,g23517);
  not NOT_9235(g24334,II31676);
  not NOT_9236(II31679,g23453);
  not NOT_9237(g24335,II31679);
  not NOT_9238(II31682,g24240);
  not NOT_9239(g24336,II31682);
  not NOT_9240(II31685,g23626);
  not NOT_9241(g24337,II31685);
  not NOT_9242(II31688,g24035);
  not NOT_9243(g24338,II31688);
  not NOT_9244(II31691,g24053);
  not NOT_9245(g24339,II31691);
  not NOT_9246(II31694,g24064);
  not NOT_9247(g24340,II31694);
  not NOT_9248(II31697,g23791);
  not NOT_9249(g24341,II31697);
  not NOT_9250(II31700,g23835);
  not NOT_9251(g24342,II31700);
  not NOT_9252(II31703,g23861);
  not NOT_9253(g24343,II31703);
  not NOT_9254(II31706,g23836);
  not NOT_9255(g24344,II31706);
  not NOT_9256(II31709,g23862);
  not NOT_9257(g24345,II31709);
  not NOT_9258(II31712,g23890);
  not NOT_9259(g24346,II31712);
  not NOT_9260(II31715,g23566);
  not NOT_9261(g24347,II31715);
  not NOT_9262(II31718,g23580);
  not NOT_9263(g24348,II31718);
  not NOT_9264(II31721,g23601);
  not NOT_9265(g24349,II31721);
  not NOT_9266(II31724,g23581);
  not NOT_9267(g24350,II31724);
  not NOT_9268(II31727,g23602);
  not NOT_9269(g24351,II31727);
  not NOT_9270(II31730,g23627);
  not NOT_9271(g24352,II31730);
  not NOT_9272(II31733,g23603);
  not NOT_9273(g24353,II31733);
  not NOT_9274(II31736,g23628);
  not NOT_9275(g24354,II31736);
  not NOT_9276(II31739,g23668);
  not NOT_9277(g24355,II31739);
  not NOT_9278(II31742,g23629);
  not NOT_9279(g24356,II31742);
  not NOT_9280(II31745,g23669);
  not NOT_9281(g24357,II31745);
  not NOT_9282(II31748,g23711);
  not NOT_9283(g24358,II31748);
  not NOT_9284(II31751,g23670);
  not NOT_9285(g24359,II31751);
  not NOT_9286(II31754,g23712);
  not NOT_9287(g24360,II31754);
  not NOT_9288(II31757,g23744);
  not NOT_9289(g24361,II31757);
  not NOT_9290(II31760,g23713);
  not NOT_9291(g24362,II31760);
  not NOT_9292(II31763,g23745);
  not NOT_9293(g24363,II31763);
  not NOT_9294(II31766,g23792);
  not NOT_9295(g24364,II31766);
  not NOT_9296(II31769,g23746);
  not NOT_9297(g24365,II31769);
  not NOT_9298(II31772,g23793);
  not NOT_9299(g24366,II31772);
  not NOT_9300(II31775,g23837);
  not NOT_9301(g24367,II31775);
  not NOT_9302(II31778,g23794);
  not NOT_9303(g24368,II31778);
  not NOT_9304(II31781,g23838);
  not NOT_9305(g24369,II31781);
  not NOT_9306(II31784,g23863);
  not NOT_9307(g24370,II31784);
  not NOT_9308(II31787,g23531);
  not NOT_9309(g24371,II31787);
  not NOT_9310(II31790,g23459);
  not NOT_9311(g24372,II31790);
  not NOT_9312(II31793,g23472);
  not NOT_9313(g24373,II31793);
  not NOT_9314(II31796,g23508);
  not NOT_9315(g24374,II31796);
  not NOT_9316(II31799,g23532);
  not NOT_9317(g24375,II31799);
  not NOT_9318(II31802,g23460);
  not NOT_9319(g24376,II31802);
  not NOT_9320(II31805,g24248);
  not NOT_9321(g24377,II31805);
  not NOT_9322(II31808,g23675);
  not NOT_9323(g24378,II31808);
  not NOT_9324(II31811,g24055);
  not NOT_9325(g24379,II31811);
  not NOT_9326(II31814,g24066);
  not NOT_9327(g24380,II31814);
  not NOT_9328(II31817,g24077);
  not NOT_9329(g24381,II31817);
  not NOT_9330(II31820,g23844);
  not NOT_9331(g24382,II31820);
  not NOT_9332(II31823,g23870);
  not NOT_9333(g24383,II31823);
  not NOT_9334(II31826,g23895);
  not NOT_9335(g24384,II31826);
  not NOT_9336(II31829,g23871);
  not NOT_9337(g24385,II31829);
  not NOT_9338(II31832,g23896);
  not NOT_9339(g24386,II31832);
  not NOT_9340(II31835,g23911);
  not NOT_9341(g24387,II31835);
  not NOT_9342(II31838,g23585);
  not NOT_9343(g24388,II31838);
  not NOT_9344(II31841,g23607);
  not NOT_9345(g24389,II31841);
  not NOT_9346(II31844,g23633);
  not NOT_9347(g24390,II31844);
  not NOT_9348(II31847,g23608);
  not NOT_9349(g24391,II31847);
  not NOT_9350(II31850,g23634);
  not NOT_9351(g24392,II31850);
  not NOT_9352(II31853,g23676);
  not NOT_9353(g24393,II31853);
  not NOT_9354(II31856,g23635);
  not NOT_9355(g24394,II31856);
  not NOT_9356(II31859,g23677);
  not NOT_9357(g24395,II31859);
  not NOT_9358(II31862,g23718);
  not NOT_9359(g24396,II31862);
  not NOT_9360(II31865,g23678);
  not NOT_9361(g24397,II31865);
  not NOT_9362(II31868,g23719);
  not NOT_9363(g24398,II31868);
  not NOT_9364(II31871,g23765);
  not NOT_9365(g24399,II31871);
  not NOT_9366(II31874,g23720);
  not NOT_9367(g24400,II31874);
  not NOT_9368(II31877,g23766);
  not NOT_9369(g24401,II31877);
  not NOT_9370(II31880,g23799);
  not NOT_9371(g24402,II31880);
  not NOT_9372(II31883,g23767);
  not NOT_9373(g24403,II31883);
  not NOT_9374(II31886,g23800);
  not NOT_9375(g24404,II31886);
  not NOT_9376(II31889,g23845);
  not NOT_9377(g24405,II31889);
  not NOT_9378(II31892,g23801);
  not NOT_9379(g24406,II31892);
  not NOT_9380(II31895,g23846);
  not NOT_9381(g24407,II31895);
  not NOT_9382(II31898,g23872);
  not NOT_9383(g24408,II31898);
  not NOT_9384(II31901,g23847);
  not NOT_9385(g24409,II31901);
  not NOT_9386(II31904,g23873);
  not NOT_9387(g24410,II31904);
  not NOT_9388(II31907,g23897);
  not NOT_9389(g24411,II31907);
  not NOT_9390(II31910,g23542);
  not NOT_9391(g24412,II31910);
  not NOT_9392(II31913,g23468);
  not NOT_9393(g24413,II31913);
  not NOT_9394(II31916,g23485);
  not NOT_9395(g24414,II31916);
  not NOT_9396(II31919,g23524);
  not NOT_9397(g24415,II31919);
  not NOT_9398(II31922,g23543);
  not NOT_9399(g24416,II31922);
  not NOT_9400(II31925,g23469);
  not NOT_9401(g24417,II31925);
  not NOT_9402(II31928,g24255);
  not NOT_9403(g24418,II31928);
  not NOT_9404(II31931,g23725);
  not NOT_9405(g24419,II31931);
  not NOT_9406(II31934,g24068);
  not NOT_9407(g24420,II31934);
  not NOT_9408(II31937,g24079);
  not NOT_9409(g24421,II31937);
  not NOT_9410(II31940,g24088);
  not NOT_9411(g24422,II31940);
  not NOT_9412(II31943,g24000);
  not NOT_9413(g24423,II31943);
  not NOT_9414(II31946,g23916);
  not NOT_9415(g24424,II31946);
  not NOT_9416(II31949,g23943);
  not NOT_9417(g24425,II31949);
  not NOT_9418(g24482,g24183);
  not NOT_9419(II32042,g23399);
  not NOT_9420(g24518,II32042);
  not NOT_9421(II32057,g23406);
  not NOT_9422(g24531,II32057);
  not NOT_9423(II32067,g24174);
  not NOT_9424(g24539,II32067);
  not NOT_9425(II32074,g23413);
  not NOT_9426(g24544,II32074);
  not NOT_9427(II32081,g24178);
  not NOT_9428(g24549,II32081);
  not NOT_9429(II32085,g24179);
  not NOT_9430(g24551,II32085);
  not NOT_9431(II32092,g23418);
  not NOT_9432(g24556,II32092);
  not NOT_9433(II32098,g24181);
  not NOT_9434(g24560,II32098);
  not NOT_9435(II32102,g24182);
  not NOT_9436(g24562,II32102);
  not NOT_9437(II32109,g24206);
  not NOT_9438(g24567,II32109);
  not NOT_9439(II32112,g24207);
  not NOT_9440(g24568,II32112);
  not NOT_9441(II32116,g24208);
  not NOT_9442(g24570,II32116);
  not NOT_9443(II32120,g24209);
  not NOT_9444(g24572,II32120);
  not NOT_9445(II32126,g24212);
  not NOT_9446(g24576,II32126);
  not NOT_9447(II32129,g24213);
  not NOT_9448(g24577,II32129);
  not NOT_9449(II32133,g24214);
  not NOT_9450(g24579,II32133);
  not NOT_9451(II32137,g24215);
  not NOT_9452(g24581,II32137);
  not NOT_9453(II32140,g24216);
  not NOT_9454(g24582,II32140);
  not NOT_9455(II32143,g24218);
  not NOT_9456(g24583,II32143);
  not NOT_9457(II32146,g24219);
  not NOT_9458(g24584,II32146);
  not NOT_9459(II32150,g24222);
  not NOT_9460(g24586,II32150);
  not NOT_9461(II32153,g24223);
  not NOT_9462(g24587,II32153);
  not NOT_9463(II32156,g24225);
  not NOT_9464(g24588,II32156);
  not NOT_9465(II32159,g24226);
  not NOT_9466(g24589,II32159);
  not NOT_9467(II32164,g24228);
  not NOT_9468(g24592,II32164);
  not NOT_9469(II32167,g24230);
  not NOT_9470(g24593,II32167);
  not NOT_9471(II32170,g24231);
  not NOT_9472(g24594,II32170);
  not NOT_9473(II32175,g24235);
  not NOT_9474(g24597,II32175);
  not NOT_9475(II32178,g24237);
  not NOT_9476(g24598,II32178);
  not NOT_9477(II32181,g24238);
  not NOT_9478(g24599,II32181);
  not NOT_9479(II32184,g23497);
  not NOT_9480(g24600,II32184);
  not NOT_9481(II32189,g24243);
  not NOT_9482(g24605,II32189);
  not NOT_9483(II32193,g23513);
  not NOT_9484(g24607,II32193);
  not NOT_9485(II32198,g24250);
  not NOT_9486(g24612,II32198);
  not NOT_9487(II32203,g23528);
  not NOT_9488(g24619,II32203);
  not NOT_9489(II32210,g23539);
  not NOT_9490(g24630,II32210);
  not NOT_9491(g24648,g23470);
  not NOT_9492(g24668,g23482);
  not NOT_9493(g24687,g23493);
  not NOT_9494(g24704,g23509);
  not NOT_9495(II32248,g23919);
  not NOT_9496(g24734,II32248);
  not NOT_9497(II32251,g23919);
  not NOT_9498(g24735,II32251);
  not NOT_9499(II32281,g23950);
  not NOT_9500(g24763,II32281);
  not NOT_9501(II32320,g23979);
  not NOT_9502(g24784,II32320);
  not NOT_9503(II32365,g24009);
  not NOT_9504(g24805,II32365);
  not NOT_9505(g24815,g23448);
  not NOT_9506(II32388,g23385);
  not NOT_9507(g24816,II32388);
  not NOT_9508(II32419,g24043);
  not NOT_9509(g24827,II32419);
  not NOT_9510(g24834,g23455);
  not NOT_9511(II32439,g23392);
  not NOT_9512(g24835,II32439);
  not NOT_9513(g24850,g23464);
  not NOT_9514(II32487,g23400);
  not NOT_9515(g24851,II32487);
  not NOT_9516(II32506,g23324);
  not NOT_9517(g24856,II32506);
  not NOT_9518(g24864,g23473);
  not NOT_9519(II32535,g23407);
  not NOT_9520(g24865,II32535);
  not NOT_9521(II32556,g23329);
  not NOT_9522(g24872,II32556);
  not NOT_9523(II32583,g23330);
  not NOT_9524(g24879,II32583);
  not NOT_9525(II32604,g23339);
  not NOT_9526(g24886,II32604);
  not NOT_9527(g24893,g23486);
  not NOT_9528(II32642,g23348);
  not NOT_9529(g24903,II32642);
  not NOT_9530(g24912,g23495);
  not NOT_9531(g24916,g23502);
  not NOT_9532(g24929,g23511);
  not NOT_9533(g24933,g23518);
  not NOT_9534(g24939,g23660);
  not NOT_9535(g24941,g23526);
  not NOT_9536(g24945,g23533);
  not NOT_9537(II32704,g23357);
  not NOT_9538(g24949,II32704);
  not NOT_9539(g24950,g23710);
  not NOT_9540(g24952,g23537);
  not NOT_9541(II32716,g23358);
  not NOT_9542(g24956,II32716);
  not NOT_9543(II32719,g23359);
  not NOT_9544(g24957,II32719);
  not NOT_9545(g24958,g23478);
  not NOT_9546(g24962,g23764);
  not NOT_9547(g24969,g23489);
  not NOT_9548(g24973,g23819);
  not NOT_9549(g24982,g23505);
  not NOT_9550(g24993,g23521);
  not NOT_9551(g25087,g23731);
  not NOT_9552(g25094,g23779);
  not NOT_9553(g25095,g23786);
  not NOT_9554(II32829,g24059);
  not NOT_9555(g25103,II32829);
  not NOT_9556(g25104,g23832);
  not NOT_9557(g25105,g23839);
  not NOT_9558(II32835,g24072);
  not NOT_9559(g25109,II32835);
  not NOT_9560(g25110,g23867);
  not NOT_9561(g25111,g23874);
  not NOT_9562(g25115,g23879);
  not NOT_9563(g25116,g23882);
  not NOT_9564(II32844,g23644);
  not NOT_9565(g25118,II32844);
  not NOT_9566(II32847,g24083);
  not NOT_9567(g25119,II32847);
  not NOT_9568(g25120,g23901);
  not NOT_9569(II32851,g23694);
  not NOT_9570(g25121,II32851);
  not NOT_9571(II32854,g24092);
  not NOT_9572(g25122,II32854);
  not NOT_9573(II32857,g23748);
  not NOT_9574(g25123,II32857);
  not NOT_9575(II32860,g23803);
  not NOT_9576(g25124,II32860);
  not NOT_9577(g25126,g24030);
  not NOT_9578(II32868,g25118);
  not NOT_9579(g25130,II32868);
  not NOT_9580(II32871,g24518);
  not NOT_9581(g25131,II32871);
  not NOT_9582(II32874,g24539);
  not NOT_9583(g25132,II32874);
  not NOT_9584(II32877,g24567);
  not NOT_9585(g25133,II32877);
  not NOT_9586(II32880,g24581);
  not NOT_9587(g25134,II32880);
  not NOT_9588(II32883,g24592);
  not NOT_9589(g25135,II32883);
  not NOT_9590(II32886,g24549);
  not NOT_9591(g25136,II32886);
  not NOT_9592(II32889,g24568);
  not NOT_9593(g25137,II32889);
  not NOT_9594(II32892,g24582);
  not NOT_9595(g25138,II32892);
  not NOT_9596(II32895,g24816);
  not NOT_9597(g25139,II32895);
  not NOT_9598(II32898,g24856);
  not NOT_9599(g25140,II32898);
  not NOT_9600(II32901,g25121);
  not NOT_9601(g25141,II32901);
  not NOT_9602(II32904,g24531);
  not NOT_9603(g25142,II32904);
  not NOT_9604(II32907,g24551);
  not NOT_9605(g25143,II32907);
  not NOT_9606(II32910,g24576);
  not NOT_9607(g25144,II32910);
  not NOT_9608(II32913,g24586);
  not NOT_9609(g25145,II32913);
  not NOT_9610(II32916,g24597);
  not NOT_9611(g25146,II32916);
  not NOT_9612(II32919,g24560);
  not NOT_9613(g25147,II32919);
  not NOT_9614(II32922,g24577);
  not NOT_9615(g25148,II32922);
  not NOT_9616(II32925,g24587);
  not NOT_9617(g25149,II32925);
  not NOT_9618(II32928,g24835);
  not NOT_9619(g25150,II32928);
  not NOT_9620(II32931,g24872);
  not NOT_9621(g25151,II32931);
  not NOT_9622(II32934,g25123);
  not NOT_9623(g25152,II32934);
  not NOT_9624(II32937,g24544);
  not NOT_9625(g25153,II32937);
  not NOT_9626(II32940,g24562);
  not NOT_9627(g25154,II32940);
  not NOT_9628(II32943,g24583);
  not NOT_9629(g25155,II32943);
  not NOT_9630(II32946,g24593);
  not NOT_9631(g25156,II32946);
  not NOT_9632(II32949,g24605);
  not NOT_9633(g25157,II32949);
  not NOT_9634(II32952,g24570);
  not NOT_9635(g25158,II32952);
  not NOT_9636(II32955,g24584);
  not NOT_9637(g25159,II32955);
  not NOT_9638(II32958,g24594);
  not NOT_9639(g25160,II32958);
  not NOT_9640(II32961,g24851);
  not NOT_9641(g25161,II32961);
  not NOT_9642(II32964,g24886);
  not NOT_9643(g25162,II32964);
  not NOT_9644(II32967,g25124);
  not NOT_9645(g25163,II32967);
  not NOT_9646(II32970,g24556);
  not NOT_9647(g25164,II32970);
  not NOT_9648(II32973,g24572);
  not NOT_9649(g25165,II32973);
  not NOT_9650(II32976,g24588);
  not NOT_9651(g25166,II32976);
  not NOT_9652(II32979,g24598);
  not NOT_9653(g25167,II32979);
  not NOT_9654(II32982,g24612);
  not NOT_9655(g25168,II32982);
  not NOT_9656(II32985,g24579);
  not NOT_9657(g25169,II32985);
  not NOT_9658(II32988,g24589);
  not NOT_9659(g25170,II32988);
  not NOT_9660(II32991,g24599);
  not NOT_9661(g25171,II32991);
  not NOT_9662(II32994,g24865);
  not NOT_9663(g25172,II32994);
  not NOT_9664(II32997,g24903);
  not NOT_9665(g25173,II32997);
  not NOT_9666(II33000,g24949);
  not NOT_9667(g25174,II33000);
  not NOT_9668(II33003,g24956);
  not NOT_9669(g25175,II33003);
  not NOT_9670(II33006,g24957);
  not NOT_9671(g25176,II33006);
  not NOT_9672(II33009,g24879);
  not NOT_9673(g25177,II33009);
  not NOT_9674(II33013,g25119);
  not NOT_9675(g25179,II33013);
  not NOT_9676(II33016,g25122);
  not NOT_9677(g25180,II33016);
  not NOT_9678(g25274,g24912);
  not NOT_9679(g25283,g24929);
  not NOT_9680(g25291,g24941);
  not NOT_9681(II33128,g24975);
  not NOT_9682(g25296,II33128);
  not NOT_9683(g25301,g24952);
  not NOT_9684(g25305,g24880);
  not NOT_9685(II33136,g24986);
  not NOT_9686(g25306,II33136);
  not NOT_9687(g25313,g24868);
  not NOT_9688(g25314,g24897);
  not NOT_9689(II33145,g24997);
  not NOT_9690(g25315,II33145);
  not NOT_9691(g25319,g24857);
  not NOT_9692(g25322,g24883);
  not NOT_9693(g25323,g24920);
  not NOT_9694(II33154,g25005);
  not NOT_9695(g25324,II33154);
  not NOT_9696(II33157,g25027);
  not NOT_9697(g25327,II33157);
  not NOT_9698(g25329,g24844);
  not NOT_9699(g25330,g24873);
  not NOT_9700(g25332,g24900);
  not NOT_9701(g25333,g24937);
  not NOT_9702(g25335,g24832);
  not NOT_9703(II33168,g25042);
  not NOT_9704(g25336,II33168);
  not NOT_9705(g25338,g24860);
  not NOT_9706(g25339,g24887);
  not NOT_9707(g25341,g24923);
  not NOT_9708(g25347,g24817);
  not NOT_9709(g25349,g24848);
  not NOT_9710(II33182,g25056);
  not NOT_9711(g25350,II33182);
  not NOT_9712(g25352,g24875);
  not NOT_9713(g25353,g24904);
  not NOT_9714(II33188,g24814);
  not NOT_9715(g25354,II33188);
  not NOT_9716(g25355,g24797);
  not NOT_9717(g25361,g24837);
  not NOT_9718(g25363,g24862);
  not NOT_9719(II33198,g25067);
  not NOT_9720(g25364,II33198);
  not NOT_9721(g25366,g24889);
  not NOT_9722(g25367,g24676);
  not NOT_9723(g25368,g24778);
  not NOT_9724(II33205,g24833);
  not NOT_9725(g25369,II33205);
  not NOT_9726(g25370,g24820);
  not NOT_9727(g25376,g24852);
  not NOT_9728(g25378,g24877);
  not NOT_9729(g25379,g24893);
  not NOT_9730(g25383,g24766);
  not NOT_9731(g25384,g24695);
  not NOT_9732(g25385,g24801);
  not NOT_9733(II33219,g24849);
  not NOT_9734(g25386,II33219);
  not NOT_9735(g25387,g24839);
  not NOT_9736(g25393,g24866);
  not NOT_9737(g25394,g24753);
  not NOT_9738(g25395,g24916);
  not NOT_9739(g25399,g24787);
  not NOT_9740(g25400,g24712);
  not NOT_9741(g25401,g24823);
  not NOT_9742(II33232,g24863);
  not NOT_9743(g25402,II33232);
  not NOT_9744(g25403,g24854);
  not NOT_9745(g25404,g24771);
  not NOT_9746(g25405,g24933);
  not NOT_9747(g25409,g24808);
  not NOT_9748(g25410,g24723);
  not NOT_9749(g25411,g24842);
  not NOT_9750(g25412,g24791);
  not NOT_9751(g25413,g24945);
  not NOT_9752(g25417,g24830);
  not NOT_9753(g25419,g24812);
  not NOT_9754(II33246,g24890);
  not NOT_9755(g25420,II33246);
  not NOT_9756(II33249,g24890);
  not NOT_9757(g25421,II33249);
  not NOT_9758(g25422,g24958);
  not NOT_9759(g25430,g24616);
  not NOT_9760(g25431,g24969);
  not NOT_9761(II33257,g24909);
  not NOT_9762(g25435,II33257);
  not NOT_9763(II33260,g24909);
  not NOT_9764(g25436,II33260);
  not NOT_9765(g25437,g24627);
  not NOT_9766(g25438,g24982);
  not NOT_9767(II33265,g24925);
  not NOT_9768(g25442,II33265);
  not NOT_9769(II33268,g24925);
  not NOT_9770(g25443,II33268);
  not NOT_9771(g25444,g24641);
  not NOT_9772(g25445,g24993);
  not NOT_9773(g25449,g24660);
  not NOT_9774(II33278,g25088);
  not NOT_9775(g25454,II33278);
  not NOT_9776(II33282,g25096);
  not NOT_9777(g25458,II33282);
  not NOT_9778(II33286,g24426);
  not NOT_9779(g25462,II33286);
  not NOT_9780(II33289,g25106);
  not NOT_9781(g25463,II33289);
  not NOT_9782(II33293,g25008);
  not NOT_9783(g25467,II33293);
  not NOT_9784(II33297,g24430);
  not NOT_9785(g25471,II33297);
  not NOT_9786(II33300,g25112);
  not NOT_9787(g25472,II33300);
  not NOT_9788(II33304,g25004);
  not NOT_9789(g25476,II33304);
  not NOT_9790(II33307,g25011);
  not NOT_9791(g25479,II33307);
  not NOT_9792(II33312,g25014);
  not NOT_9793(g25484,II33312);
  not NOT_9794(II33316,g24434);
  not NOT_9795(g25488,II33316);
  not NOT_9796(II33321,g24442);
  not NOT_9797(g25493,II33321);
  not NOT_9798(II33324,g25009);
  not NOT_9799(g25496,II33324);
  not NOT_9800(II33327,g25017);
  not NOT_9801(g25499,II33327);
  not NOT_9802(II33330,g25019);
  not NOT_9803(g25502,II33330);
  not NOT_9804(II33335,g25010);
  not NOT_9805(g25507,II33335);
  not NOT_9806(II33338,g25021);
  not NOT_9807(g25510,II33338);
  not NOT_9808(II33343,g25024);
  not NOT_9809(g25515,II33343);
  not NOT_9810(II33347,g24438);
  not NOT_9811(g25519,II33347);
  not NOT_9812(II33352,g24443);
  not NOT_9813(g25524,II33352);
  not NOT_9814(II33355,g25012);
  not NOT_9815(g25527,II33355);
  not NOT_9816(II33358,g25028);
  not NOT_9817(g25530,II33358);
  not NOT_9818(II33361,g25013);
  not NOT_9819(g25533,II33361);
  not NOT_9820(II33364,g25029);
  not NOT_9821(g25536,II33364);
  not NOT_9822(II33368,g24444);
  not NOT_9823(g25540,II33368);
  not NOT_9824(II33371,g25015);
  not NOT_9825(g25543,II33371);
  not NOT_9826(II33374,g25031);
  not NOT_9827(g25546,II33374);
  not NOT_9828(II33377,g25033);
  not NOT_9829(g25549,II33377);
  not NOT_9830(II33382,g25016);
  not NOT_9831(g25554,II33382);
  not NOT_9832(II33385,g25035);
  not NOT_9833(g25557,II33385);
  not NOT_9834(II33390,g25038);
  not NOT_9835(g25562,II33390);
  not NOT_9836(II33396,g24447);
  not NOT_9837(g25573,II33396);
  not NOT_9838(II33399,g25018);
  not NOT_9839(g25576,II33399);
  not NOT_9840(II33402,g24448);
  not NOT_9841(g25579,II33402);
  not NOT_9842(II33405,g25020);
  not NOT_9843(g25582,II33405);
  not NOT_9844(II33408,g25040);
  not NOT_9845(g25585,II33408);
  not NOT_9846(II33411,g24491);
  not NOT_9847(g25588,II33411);
  not NOT_9848(II33415,g24449);
  not NOT_9849(g25590,II33415);
  not NOT_9850(II33418,g25022);
  not NOT_9851(g25593,II33418);
  not NOT_9852(II33421,g25043);
  not NOT_9853(g25596,II33421);
  not NOT_9854(II33424,g25023);
  not NOT_9855(g25599,II33424);
  not NOT_9856(II33427,g25044);
  not NOT_9857(g25602,II33427);
  not NOT_9858(II33431,g24450);
  not NOT_9859(g25606,II33431);
  not NOT_9860(II33434,g25025);
  not NOT_9861(g25609,II33434);
  not NOT_9862(II33437,g25046);
  not NOT_9863(g25612,II33437);
  not NOT_9864(II33440,g25048);
  not NOT_9865(g25615,II33440);
  not NOT_9866(II33445,g25026);
  not NOT_9867(g25620,II33445);
  not NOT_9868(II33448,g25050);
  not NOT_9869(g25623,II33448);
  not NOT_9870(g25630,g24478);
  not NOT_9871(II33457,g24451);
  not NOT_9872(g25634,II33457);
  not NOT_9873(II33460,g24452);
  not NOT_9874(g25637,II33460);
  not NOT_9875(II33463,g25030);
  not NOT_9876(g25640,II33463);
  not NOT_9877(II33466,g25053);
  not NOT_9878(g25643,II33466);
  not NOT_9879(II33469,g24498);
  not NOT_9880(g25646,II33469);
  not NOT_9881(II33472,g24499);
  not NOT_9882(g25647,II33472);
  not NOT_9883(II33476,g24453);
  not NOT_9884(g25652,II33476);
  not NOT_9885(II33479,g25032);
  not NOT_9886(g25655,II33479);
  not NOT_9887(II33482,g24454);
  not NOT_9888(g25658,II33482);
  not NOT_9889(II33485,g25034);
  not NOT_9890(g25661,II33485);
  not NOT_9891(II33488,g25054);
  not NOT_9892(g25664,II33488);
  not NOT_9893(II33491,g24501);
  not NOT_9894(g25667,II33491);
  not NOT_9895(II33495,g24455);
  not NOT_9896(g25669,II33495);
  not NOT_9897(II33498,g25036);
  not NOT_9898(g25672,II33498);
  not NOT_9899(II33501,g25057);
  not NOT_9900(g25675,II33501);
  not NOT_9901(II33504,g25037);
  not NOT_9902(g25678,II33504);
  not NOT_9903(II33507,g25058);
  not NOT_9904(g25681,II33507);
  not NOT_9905(II33511,g24456);
  not NOT_9906(g25685,II33511);
  not NOT_9907(II33514,g25039);
  not NOT_9908(g25688,II33514);
  not NOT_9909(II33517,g25060);
  not NOT_9910(g25691,II33517);
  not NOT_9911(II33520,g25062);
  not NOT_9912(g25694,II33520);
  not NOT_9913(g25698,g24600);
  not NOT_9914(II33526,g24457);
  not NOT_9915(g25700,II33526);
  not NOT_9916(II33529,g25041);
  not NOT_9917(g25703,II33529);
  not NOT_9918(II33532,g24507);
  not NOT_9919(g25706,II33532);
  not NOT_9920(II33535,g24508);
  not NOT_9921(g25707,II33535);
  not NOT_9922(II33539,g24458);
  not NOT_9923(g25711,II33539);
  not NOT_9924(II33542,g24459);
  not NOT_9925(g25714,II33542);
  not NOT_9926(II33545,g25045);
  not NOT_9927(g25717,II33545);
  not NOT_9928(II33548,g25064);
  not NOT_9929(g25720,II33548);
  not NOT_9930(II33551,g24510);
  not NOT_9931(g25723,II33551);
  not NOT_9932(II33554,g24511);
  not NOT_9933(g25724,II33554);
  not NOT_9934(II33558,g24460);
  not NOT_9935(g25729,II33558);
  not NOT_9936(II33561,g25047);
  not NOT_9937(g25732,II33561);
  not NOT_9938(II33564,g24461);
  not NOT_9939(g25735,II33564);
  not NOT_9940(II33567,g25049);
  not NOT_9941(g25738,II33567);
  not NOT_9942(II33570,g25065);
  not NOT_9943(g25741,II33570);
  not NOT_9944(II33573,g24513);
  not NOT_9945(g25744,II33573);
  not NOT_9946(II33577,g24462);
  not NOT_9947(g25746,II33577);
  not NOT_9948(II33580,g25051);
  not NOT_9949(g25749,II33580);
  not NOT_9950(II33583,g25068);
  not NOT_9951(g25752,II33583);
  not NOT_9952(II33586,g25052);
  not NOT_9953(g25755,II33586);
  not NOT_9954(II33589,g25069);
  not NOT_9955(g25758,II33589);
  not NOT_9956(II33593,g24445);
  not NOT_9957(g25762,II33593);
  not NOT_9958(II33596,g24446);
  not NOT_9959(g25763,II33596);
  not NOT_9960(II33600,g24463);
  not NOT_9961(g25767,II33600);
  not NOT_9962(II33603,g24519);
  not NOT_9963(g25770,II33603);
  not NOT_9964(g25771,g24607);
  not NOT_9965(II33608,g24464);
  not NOT_9966(g25773,II33608);
  not NOT_9967(II33611,g25055);
  not NOT_9968(g25776,II33611);
  not NOT_9969(II33614,g24521);
  not NOT_9970(g25779,II33614);
  not NOT_9971(II33617,g24522);
  not NOT_9972(g25780,II33617);
  not NOT_9973(II33621,g24465);
  not NOT_9974(g25784,II33621);
  not NOT_9975(II33624,g24466);
  not NOT_9976(g25787,II33624);
  not NOT_9977(II33627,g25059);
  not NOT_9978(g25790,II33627);
  not NOT_9979(II33630,g25071);
  not NOT_9980(g25793,II33630);
  not NOT_9981(II33633,g24524);
  not NOT_9982(g25796,II33633);
  not NOT_9983(II33636,g24525);
  not NOT_9984(g25797,II33636);
  not NOT_9985(II33640,g24467);
  not NOT_9986(g25802,II33640);
  not NOT_9987(II33643,g25061);
  not NOT_9988(g25805,II33643);
  not NOT_9989(II33646,g24468);
  not NOT_9990(g25808,II33646);
  not NOT_9991(II33649,g25063);
  not NOT_9992(g25811,II33649);
  not NOT_9993(II33652,g25072);
  not NOT_9994(g25814,II33652);
  not NOT_9995(II33655,g24527);
  not NOT_9996(g25817,II33655);
  not NOT_9997(II33659,g24469);
  not NOT_9998(g25821,II33659);
  not NOT_9999(II33662,g24532);
  not NOT_10000(g25824,II33662);
  not NOT_10001(g25825,g24619);
  not NOT_10002(II33667,g24470);
  not NOT_10003(g25827,II33667);
  not NOT_10004(II33670,g25066);
  not NOT_10005(g25830,II33670);
  not NOT_10006(II33673,g24534);
  not NOT_10007(g25833,II33673);
  not NOT_10008(II33676,g24535);
  not NOT_10009(g25834,II33676);
  not NOT_10010(II33680,g24471);
  not NOT_10011(g25838,II33680);
  not NOT_10012(II33683,g24472);
  not NOT_10013(g25841,II33683);
  not NOT_10014(II33686,g25070);
  not NOT_10015(g25844,II33686);
  not NOT_10016(II33689,g25074);
  not NOT_10017(g25847,II33689);
  not NOT_10018(II33692,g24537);
  not NOT_10019(g25850,II33692);
  not NOT_10020(II33695,g24538);
  not NOT_10021(g25851,II33695);
  not NOT_10022(II33700,g24474);
  not NOT_10023(g25856,II33700);
  not NOT_10024(II33703,g24545);
  not NOT_10025(g25859,II33703);
  not NOT_10026(g25860,g24630);
  not NOT_10027(II33708,g24475);
  not NOT_10028(g25862,II33708);
  not NOT_10029(II33711,g25073);
  not NOT_10030(g25865,II33711);
  not NOT_10031(II33714,g24547);
  not NOT_10032(g25868,II33714);
  not NOT_10033(II33717,g24548);
  not NOT_10034(g25869,II33717);
  not NOT_10035(II33723,g24477);
  not NOT_10036(g25877,II33723);
  not NOT_10037(II33726,g24557);
  not NOT_10038(g25880,II33726);
  not NOT_10039(II33732,g24473);
  not NOT_10040(g25886,II33732);
  not NOT_10041(II33737,g24476);
  not NOT_10042(g25891,II33737);
  not NOT_10043(g25895,g24939);
  not NOT_10044(g25899,g24928);
  not NOT_10045(g25903,g24950);
  not NOT_10046(g25907,g24940);
  not NOT_10047(g25911,g24962);
  not NOT_10048(g25915,g24951);
  not NOT_10049(g25919,g24973);
  not NOT_10050(g25923,g24963);
  not NOT_10051(g25937,g24763);
  not NOT_10052(g25939,g24784);
  not NOT_10053(g25942,g24805);
  not NOT_10054(g25945,g24827);
  not NOT_10055(g25952,g24735);
  not NOT_10056(II33790,g25103);
  not NOT_10057(g25976,II33790);
  not NOT_10058(II33798,g25109);
  not NOT_10059(g25982,II33798);
  not NOT_10060(II33801,g25327);
  not NOT_10061(g25983,II33801);
  not NOT_10062(II33804,g25976);
  not NOT_10063(g25984,II33804);
  not NOT_10064(II33807,g25588);
  not NOT_10065(g25985,II33807);
  not NOT_10066(II33810,g25646);
  not NOT_10067(g25986,II33810);
  not NOT_10068(II33813,g25706);
  not NOT_10069(g25987,II33813);
  not NOT_10070(II33816,g25647);
  not NOT_10071(g25988,II33816);
  not NOT_10072(II33819,g25707);
  not NOT_10073(g25989,II33819);
  not NOT_10074(II33822,g25770);
  not NOT_10075(g25990,II33822);
  not NOT_10076(II33825,g25462);
  not NOT_10077(g25991,II33825);
  not NOT_10078(II33828,g25336);
  not NOT_10079(g25992,II33828);
  not NOT_10080(II33831,g25982);
  not NOT_10081(g25993,II33831);
  not NOT_10082(II33834,g25667);
  not NOT_10083(g25994,II33834);
  not NOT_10084(II33837,g25723);
  not NOT_10085(g25995,II33837);
  not NOT_10086(II33840,g25779);
  not NOT_10087(g25996,II33840);
  not NOT_10088(II33843,g25724);
  not NOT_10089(g25997,II33843);
  not NOT_10090(II33846,g25780);
  not NOT_10091(g25998,II33846);
  not NOT_10092(II33849,g25824);
  not NOT_10093(g25999,II33849);
  not NOT_10094(II33852,g25471);
  not NOT_10095(g26000,II33852);
  not NOT_10096(II33855,g25350);
  not NOT_10097(g26001,II33855);
  not NOT_10098(II33858,g25179);
  not NOT_10099(g26002,II33858);
  not NOT_10100(II33861,g25744);
  not NOT_10101(g26003,II33861);
  not NOT_10102(II33864,g25796);
  not NOT_10103(g26004,II33864);
  not NOT_10104(II33867,g25833);
  not NOT_10105(g26005,II33867);
  not NOT_10106(II33870,g25797);
  not NOT_10107(g26006,II33870);
  not NOT_10108(II33873,g25834);
  not NOT_10109(g26007,II33873);
  not NOT_10110(II33876,g25859);
  not NOT_10111(g26008,II33876);
  not NOT_10112(II33879,g25488);
  not NOT_10113(g26009,II33879);
  not NOT_10114(II33882,g25364);
  not NOT_10115(g26010,II33882);
  not NOT_10116(II33885,g25180);
  not NOT_10117(g26011,II33885);
  not NOT_10118(II33888,g25817);
  not NOT_10119(g26012,II33888);
  not NOT_10120(II33891,g25850);
  not NOT_10121(g26013,II33891);
  not NOT_10122(II33894,g25868);
  not NOT_10123(g26014,II33894);
  not NOT_10124(II33897,g25851);
  not NOT_10125(g26015,II33897);
  not NOT_10126(II33900,g25869);
  not NOT_10127(g26016,II33900);
  not NOT_10128(II33903,g25880);
  not NOT_10129(g26017,II33903);
  not NOT_10130(II33906,g25519);
  not NOT_10131(g26018,II33906);
  not NOT_10132(II33909,g25886);
  not NOT_10133(g26019,II33909);
  not NOT_10134(II33912,g25891);
  not NOT_10135(g26020,II33912);
  not NOT_10136(II33915,g25762);
  not NOT_10137(g26021,II33915);
  not NOT_10138(II33918,g25763);
  not NOT_10139(g26022,II33918);
  not NOT_10140(II33954,g25343);
  not NOT_10141(g26056,II33954);
  not NOT_10142(II33961,g25357);
  not NOT_10143(g26063,II33961);
  not NOT_10144(II33968,g25372);
  not NOT_10145(g26070,II33968);
  not NOT_10146(II33974,g25389);
  not NOT_10147(g26076,II33974);
  not NOT_10148(II33984,g25932);
  not NOT_10149(g26086,II33984);
  not NOT_10150(II33990,g25870);
  not NOT_10151(g26092,II33990);
  not NOT_10152(II33995,g25935);
  not NOT_10153(g26102,II33995);
  not NOT_10154(II33999,g25490);
  not NOT_10155(g26104,II33999);
  not NOT_10156(II34002,g25490);
  not NOT_10157(g26105,II34002);
  not NOT_10158(II34009,g25882);
  not NOT_10159(g26114,II34009);
  not NOT_10160(II34012,g25938);
  not NOT_10161(g26118,II34012);
  not NOT_10162(II34017,g25887);
  not NOT_10163(g26121,II34017);
  not NOT_10164(II34020,g25940);
  not NOT_10165(g26125,II34020);
  not NOT_10166(II34026,g25892);
  not NOT_10167(g26131,II34026);
  not NOT_10168(II34029,g25520);
  not NOT_10169(g26135,II34029);
  not NOT_10170(II34032,g25520);
  not NOT_10171(g26136,II34032);
  not NOT_10172(II34041,g25566);
  not NOT_10173(g26149,II34041);
  not NOT_10174(II34044,g25566);
  not NOT_10175(g26150,II34044);
  not NOT_10176(II34051,g25204);
  not NOT_10177(g26159,II34051);
  not NOT_10178(II34056,g25206);
  not NOT_10179(g26164,II34056);
  not NOT_10180(II34059,g25207);
  not NOT_10181(g26165,II34059);
  not NOT_10182(II34063,g25209);
  not NOT_10183(g26167,II34063);
  not NOT_10184(II34068,g25211);
  not NOT_10185(g26172,II34068);
  not NOT_10186(II34071,g25212);
  not NOT_10187(g26173,II34071);
  not NOT_10188(II34074,g25213);
  not NOT_10189(g26174,II34074);
  not NOT_10190(II34077,g25954);
  not NOT_10191(g26175,II34077);
  not NOT_10192(II34080,g25539);
  not NOT_10193(g26178,II34080);
  not NOT_10194(II34083,g25214);
  not NOT_10195(g26181,II34083);
  not NOT_10196(II34086,g25215);
  not NOT_10197(g26182,II34086);
  not NOT_10198(II34091,g25217);
  not NOT_10199(g26187,II34091);
  not NOT_10200(g26189,g25952);
  not NOT_10201(II34096,g25218);
  not NOT_10202(g26190,II34096);
  not NOT_10203(II34099,g25219);
  not NOT_10204(g26191,II34099);
  not NOT_10205(II34102,g25220);
  not NOT_10206(g26192,II34102);
  not NOT_10207(II34105,g25221);
  not NOT_10208(g26193,II34105);
  not NOT_10209(II34108,g25222);
  not NOT_10210(g26194,II34108);
  not NOT_10211(II34111,g25223);
  not NOT_10212(g26195,II34111);
  not NOT_10213(II34114,g25958);
  not NOT_10214(g26196,II34114);
  not NOT_10215(II34118,g25605);
  not NOT_10216(g26202,II34118);
  not NOT_10217(II34121,g25224);
  not NOT_10218(g26205,II34121);
  not NOT_10219(II34124,g25225);
  not NOT_10220(g26206,II34124);
  not NOT_10221(II34128,g25227);
  not NOT_10222(g26208,II34128);
  not NOT_10223(g26209,g25296);
  not NOT_10224(II34132,g25228);
  not NOT_10225(g26210,II34132);
  not NOT_10226(II34135,g25229);
  not NOT_10227(g26211,II34135);
  not NOT_10228(II34140,g25230);
  not NOT_10229(g26214,II34140);
  not NOT_10230(II34143,g25231);
  not NOT_10231(g26215,II34143);
  not NOT_10232(II34146,g25232);
  not NOT_10233(g26216,II34146);
  not NOT_10234(II34150,g25233);
  not NOT_10235(g26220,II34150);
  not NOT_10236(II34153,g25234);
  not NOT_10237(g26221,II34153);
  not NOT_10238(II34156,g25235);
  not NOT_10239(g26222,II34156);
  not NOT_10240(II34159,g25964);
  not NOT_10241(g26223,II34159);
  not NOT_10242(II34162,g25684);
  not NOT_10243(g26226,II34162);
  not NOT_10244(II34165,g25236);
  not NOT_10245(g26229,II34165);
  not NOT_10246(II34168,g25237);
  not NOT_10247(g26230,II34168);
  not NOT_10248(II34172,g25239);
  not NOT_10249(g26232,II34172);
  not NOT_10250(g26237,g25306);
  not NOT_10251(II34180,g25240);
  not NOT_10252(g26238,II34180);
  not NOT_10253(II34183,g25241);
  not NOT_10254(g26239,II34183);
  not NOT_10255(II34189,g25242);
  not NOT_10256(g26245,II34189);
  not NOT_10257(II34192,g25243);
  not NOT_10258(g26246,II34192);
  not NOT_10259(II34195,g25244);
  not NOT_10260(g26247,II34195);
  not NOT_10261(II34198,g25245);
  not NOT_10262(g26248,II34198);
  not NOT_10263(II34201,g25246);
  not NOT_10264(g26249,II34201);
  not NOT_10265(II34204,g25247);
  not NOT_10266(g26250,II34204);
  not NOT_10267(II34207,g25969);
  not NOT_10268(g26251,II34207);
  not NOT_10269(II34210,g25761);
  not NOT_10270(g26254,II34210);
  not NOT_10271(II34220,g25248);
  not NOT_10272(g26264,II34220);
  not NOT_10273(g26275,g25315);
  not NOT_10274(II34230,g25249);
  not NOT_10275(g26276,II34230);
  not NOT_10276(II34233,g25250);
  not NOT_10277(g26277,II34233);
  not NOT_10278(II34238,g25251);
  not NOT_10279(g26280,II34238);
  not NOT_10280(II34241,g25252);
  not NOT_10281(g26281,II34241);
  not NOT_10282(II34244,g25253);
  not NOT_10283(g26282,II34244);
  not NOT_10284(II34254,g25185);
  not NOT_10285(g26294,II34254);
  not NOT_10286(II34266,g25255);
  not NOT_10287(g26308,II34266);
  not NOT_10288(g26313,g25324);
  not NOT_10289(II34274,g25256);
  not NOT_10290(g26314,II34274);
  not NOT_10291(II34277,g25257);
  not NOT_10292(g26315,II34277);
  not NOT_10293(II34296,g25189);
  not NOT_10294(g26341,II34296);
  not NOT_10295(II34306,g25259);
  not NOT_10296(g26349,II34306);
  not NOT_10297(II34313,g25265);
  not NOT_10298(g26354,II34313);
  not NOT_10299(II34316,g25191);
  not NOT_10300(g26355,II34316);
  not NOT_10301(II34321,g25928);
  not NOT_10302(g26358,II34321);
  not NOT_10303(II34327,g25260);
  not NOT_10304(g26364,II34327);
  not NOT_10305(II34343,g25194);
  not NOT_10306(g26385,II34343);
  not NOT_10307(II34353,g25927);
  not NOT_10308(g26393,II34353);
  not NOT_10309(II34358,g25262);
  not NOT_10310(g26398,II34358);
  not NOT_10311(II34363,g25930);
  not NOT_10312(g26401,II34363);
  not NOT_10313(II34369,g25263);
  not NOT_10314(g26407,II34369);
  not NOT_10315(II34385,g25197);
  not NOT_10316(g26428,II34385);
  not NOT_10317(II34388,g25200);
  not NOT_10318(g26429,II34388);
  not NOT_10319(II34392,g25266);
  not NOT_10320(g26433,II34392);
  not NOT_10321(II34395,g25929);
  not NOT_10322(g26434,II34395);
  not NOT_10323(II34400,g25267);
  not NOT_10324(g26439,II34400);
  not NOT_10325(II34405,g25933);
  not NOT_10326(g26442,II34405);
  not NOT_10327(II34411,g25268);
  not NOT_10328(g26448,II34411);
  not NOT_10329(II34421,g25203);
  not NOT_10330(g26461,II34421);
  not NOT_10331(II34425,g25270);
  not NOT_10332(g26465,II34425);
  not NOT_10333(II34428,g25931);
  not NOT_10334(g26466,II34428);
  not NOT_10335(II34433,g25271);
  not NOT_10336(g26471,II34433);
  not NOT_10337(II34438,g25936);
  not NOT_10338(g26474,II34438);
  not NOT_10339(II34444,g25272);
  not NOT_10340(g26480,II34444);
  not NOT_10341(g26481,g25764);
  not NOT_10342(II34449,g25205);
  not NOT_10343(g26485,II34449);
  not NOT_10344(II34453,g25279);
  not NOT_10345(g26489,II34453);
  not NOT_10346(II34456,g25934);
  not NOT_10347(g26490,II34456);
  not NOT_10348(II34461,g25280);
  not NOT_10349(g26495,II34461);
  not NOT_10350(II34464,g25199);
  not NOT_10351(g26496,II34464);
  not NOT_10352(g26497,g25818);
  not NOT_10353(II34469,g25210);
  not NOT_10354(g26501,II34469);
  not NOT_10355(II34473,g25288);
  not NOT_10356(g26505,II34473);
  not NOT_10357(II34476,g25201);
  not NOT_10358(g26506,II34476);
  not NOT_10359(II34479,g25202);
  not NOT_10360(g26507,II34479);
  not NOT_10361(g26508,g25312);
  not NOT_10362(g26512,g25853);
  not NOT_10363(g26516,g25320);
  not NOT_10364(g26520,g25874);
  not NOT_10365(g26521,g25331);
  not NOT_10366(g26525,g25340);
  not NOT_10367(g26533,g25454);
  not NOT_10368(g26538,g25458);
  not NOT_10369(g26539,g25463);
  not NOT_10370(g26540,g25467);
  not NOT_10371(g26542,g25472);
  not NOT_10372(g26543,g25476);
  not NOT_10373(g26544,g25479);
  not NOT_10374(g26546,g25484);
  not NOT_10375(II34505,g25450);
  not NOT_10376(g26548,II34505);
  not NOT_10377(g26549,g25421);
  not NOT_10378(g26550,g25493);
  not NOT_10379(g26551,g25496);
  not NOT_10380(g26552,g25499);
  not NOT_10381(g26554,g25502);
  not NOT_10382(g26555,g25507);
  not NOT_10383(g26556,g25510);
  not NOT_10384(g26558,g25515);
  not NOT_10385(g26561,g25524);
  not NOT_10386(g26562,g25527);
  not NOT_10387(g26563,g25530);
  not NOT_10388(g26564,g25533);
  not NOT_10389(g26565,g25536);
  not NOT_10390(g26566,g25540);
  not NOT_10391(g26567,g25543);
  not NOT_10392(g26568,g25546);
  not NOT_10393(g26570,g25549);
  not NOT_10394(g26571,g25554);
  not NOT_10395(g26572,g25557);
  not NOT_10396(g26574,g25562);
  not NOT_10397(II34535,g25451);
  not NOT_10398(g26576,II34535);
  not NOT_10399(g26577,g25436);
  not NOT_10400(g26578,g25573);
  not NOT_10401(g26579,g25576);
  not NOT_10402(g26580,g25579);
  not NOT_10403(g26581,g25582);
  not NOT_10404(g26582,g25585);
  not NOT_10405(g26584,g25590);
  not NOT_10406(g26585,g25593);
  not NOT_10407(g26586,g25596);
  not NOT_10408(g26587,g25599);
  not NOT_10409(g26588,g25602);
  not NOT_10410(g26589,g25606);
  not NOT_10411(g26590,g25609);
  not NOT_10412(g26591,g25612);
  not NOT_10413(g26593,g25615);
  not NOT_10414(g26594,g25620);
  not NOT_10415(g26595,g25623);
  not NOT_10416(g26597,g25443);
  not NOT_10417(g26598,g25634);
  not NOT_10418(g26599,g25637);
  not NOT_10419(g26600,g25640);
  not NOT_10420(g26601,g25643);
  not NOT_10421(g26602,g25652);
  not NOT_10422(g26603,g25655);
  not NOT_10423(g26604,g25658);
  not NOT_10424(g26605,g25661);
  not NOT_10425(g26606,g25664);
  not NOT_10426(g26608,g25669);
  not NOT_10427(g26609,g25672);
  not NOT_10428(g26610,g25675);
  not NOT_10429(g26611,g25678);
  not NOT_10430(g26612,g25681);
  not NOT_10431(g26613,g25685);
  not NOT_10432(g26614,g25688);
  not NOT_10433(g26615,g25691);
  not NOT_10434(g26617,g25694);
  not NOT_10435(II34579,g25452);
  not NOT_10436(g26618,II34579);
  not NOT_10437(g26619,g25700);
  not NOT_10438(g26620,g25703);
  not NOT_10439(g26621,g25711);
  not NOT_10440(g26622,g25714);
  not NOT_10441(g26623,g25717);
  not NOT_10442(g26624,g25720);
  not NOT_10443(g26625,g25729);
  not NOT_10444(g26626,g25732);
  not NOT_10445(g26627,g25735);
  not NOT_10446(g26628,g25738);
  not NOT_10447(g26629,g25741);
  not NOT_10448(g26631,g25746);
  not NOT_10449(g26632,g25749);
  not NOT_10450(g26633,g25752);
  not NOT_10451(g26634,g25755);
  not NOT_10452(g26635,g25758);
  not NOT_10453(g26636,g25767);
  not NOT_10454(g26637,g25773);
  not NOT_10455(g26638,g25776);
  not NOT_10456(g26639,g25784);
  not NOT_10457(g26640,g25787);
  not NOT_10458(g26641,g25790);
  not NOT_10459(g26642,g25793);
  not NOT_10460(g26643,g25802);
  not NOT_10461(g26644,g25805);
  not NOT_10462(g26645,g25808);
  not NOT_10463(g26646,g25811);
  not NOT_10464(g26647,g25814);
  not NOT_10465(g26648,g25821);
  not NOT_10466(g26649,g25827);
  not NOT_10467(g26650,g25830);
  not NOT_10468(g26651,g25838);
  not NOT_10469(g26652,g25841);
  not NOT_10470(g26653,g25844);
  not NOT_10471(g26654,g25847);
  not NOT_10472(g26656,g25856);
  not NOT_10473(g26657,g25862);
  not NOT_10474(g26658,g25865);
  not NOT_10475(g26662,g25877);
  not NOT_10476(II34641,g26086);
  not NOT_10477(g26678,II34641);
  not NOT_10478(II34644,g26159);
  not NOT_10479(g26679,II34644);
  not NOT_10480(II34647,g26164);
  not NOT_10481(g26680,II34647);
  not NOT_10482(II34650,g26172);
  not NOT_10483(g26681,II34650);
  not NOT_10484(II34653,g26165);
  not NOT_10485(g26682,II34653);
  not NOT_10486(II34656,g26173);
  not NOT_10487(g26683,II34656);
  not NOT_10488(II34659,g26190);
  not NOT_10489(g26684,II34659);
  not NOT_10490(II34662,g26174);
  not NOT_10491(g26685,II34662);
  not NOT_10492(II34665,g26191);
  not NOT_10493(g26686,II34665);
  not NOT_10494(II34668,g26210);
  not NOT_10495(g26687,II34668);
  not NOT_10496(II34671,g26192);
  not NOT_10497(g26688,II34671);
  not NOT_10498(II34674,g26211);
  not NOT_10499(g26689,II34674);
  not NOT_10500(II34677,g26232);
  not NOT_10501(g26690,II34677);
  not NOT_10502(II34680,g26294);
  not NOT_10503(g26691,II34680);
  not NOT_10504(II34683,g26364);
  not NOT_10505(g26692,II34683);
  not NOT_10506(II34686,g26398);
  not NOT_10507(g26693,II34686);
  not NOT_10508(II34689,g26433);
  not NOT_10509(g26694,II34689);
  not NOT_10510(II34692,g26102);
  not NOT_10511(g26695,II34692);
  not NOT_10512(II34695,g26167);
  not NOT_10513(g26696,II34695);
  not NOT_10514(II34698,g26181);
  not NOT_10515(g26697,II34698);
  not NOT_10516(II34701,g26193);
  not NOT_10517(g26698,II34701);
  not NOT_10518(II34704,g26182);
  not NOT_10519(g26699,II34704);
  not NOT_10520(II34707,g26194);
  not NOT_10521(g26700,II34707);
  not NOT_10522(II34710,g26214);
  not NOT_10523(g26701,II34710);
  not NOT_10524(II34713,g26195);
  not NOT_10525(g26702,II34713);
  not NOT_10526(II34716,g26215);
  not NOT_10527(g26703,II34716);
  not NOT_10528(II34719,g26238);
  not NOT_10529(g26704,II34719);
  not NOT_10530(II34722,g26216);
  not NOT_10531(g26705,II34722);
  not NOT_10532(II34725,g26239);
  not NOT_10533(g26706,II34725);
  not NOT_10534(II34728,g26264);
  not NOT_10535(g26707,II34728);
  not NOT_10536(II34731,g26341);
  not NOT_10537(g26708,II34731);
  not NOT_10538(II34734,g26407);
  not NOT_10539(g26709,II34734);
  not NOT_10540(II34737,g26439);
  not NOT_10541(g26710,II34737);
  not NOT_10542(II34740,g26465);
  not NOT_10543(g26711,II34740);
  not NOT_10544(II34743,g26118);
  not NOT_10545(g26712,II34743);
  not NOT_10546(II34746,g26187);
  not NOT_10547(g26713,II34746);
  not NOT_10548(II34749,g26205);
  not NOT_10549(g26714,II34749);
  not NOT_10550(II34752,g26220);
  not NOT_10551(g26715,II34752);
  not NOT_10552(II34755,g26206);
  not NOT_10553(g26716,II34755);
  not NOT_10554(II34758,g26221);
  not NOT_10555(g26717,II34758);
  not NOT_10556(II34761,g26245);
  not NOT_10557(g26718,II34761);
  not NOT_10558(II34764,g26222);
  not NOT_10559(g26719,II34764);
  not NOT_10560(II34767,g26246);
  not NOT_10561(g26720,II34767);
  not NOT_10562(II34770,g26276);
  not NOT_10563(g26721,II34770);
  not NOT_10564(II34773,g26247);
  not NOT_10565(g26722,II34773);
  not NOT_10566(II34776,g26277);
  not NOT_10567(g26723,II34776);
  not NOT_10568(II34779,g26308);
  not NOT_10569(g26724,II34779);
  not NOT_10570(II34782,g26385);
  not NOT_10571(g26725,II34782);
  not NOT_10572(II34785,g26448);
  not NOT_10573(g26726,II34785);
  not NOT_10574(II34788,g26471);
  not NOT_10575(g26727,II34788);
  not NOT_10576(II34791,g26489);
  not NOT_10577(g26728,II34791);
  not NOT_10578(II34794,g26125);
  not NOT_10579(g26729,II34794);
  not NOT_10580(II34797,g26208);
  not NOT_10581(g26730,II34797);
  not NOT_10582(II34800,g26229);
  not NOT_10583(g26731,II34800);
  not NOT_10584(II34803,g26248);
  not NOT_10585(g26732,II34803);
  not NOT_10586(II34806,g26230);
  not NOT_10587(g26733,II34806);
  not NOT_10588(II34809,g26249);
  not NOT_10589(g26734,II34809);
  not NOT_10590(II34812,g26280);
  not NOT_10591(g26735,II34812);
  not NOT_10592(II34815,g26250);
  not NOT_10593(g26736,II34815);
  not NOT_10594(II34818,g26281);
  not NOT_10595(g26737,II34818);
  not NOT_10596(II34821,g26314);
  not NOT_10597(g26738,II34821);
  not NOT_10598(II34824,g26282);
  not NOT_10599(g26739,II34824);
  not NOT_10600(II34827,g26315);
  not NOT_10601(g26740,II34827);
  not NOT_10602(II34830,g26349);
  not NOT_10603(g26741,II34830);
  not NOT_10604(II34833,g26428);
  not NOT_10605(g26742,II34833);
  not NOT_10606(II34836,g26480);
  not NOT_10607(g26743,II34836);
  not NOT_10608(II34839,g26495);
  not NOT_10609(g26744,II34839);
  not NOT_10610(II34842,g26505);
  not NOT_10611(g26745,II34842);
  not NOT_10612(II34845,g26496);
  not NOT_10613(g26746,II34845);
  not NOT_10614(II34848,g26506);
  not NOT_10615(g26747,II34848);
  not NOT_10616(II34851,g26354);
  not NOT_10617(g26748,II34851);
  not NOT_10618(II34854,g26507);
  not NOT_10619(g26749,II34854);
  not NOT_10620(II34857,g26355);
  not NOT_10621(g26750,II34857);
  not NOT_10622(II34860,g26548);
  not NOT_10623(g26751,II34860);
  not NOT_10624(II34863,g26576);
  not NOT_10625(g26752,II34863);
  not NOT_10626(II34866,g26618);
  not NOT_10627(g26753,II34866);
  not NOT_10628(II34872,g26217);
  not NOT_10629(g26757,II34872);
  not NOT_10630(II34879,g26240);
  not NOT_10631(g26762,II34879);
  not NOT_10632(II34901,g26295);
  not NOT_10633(g26782,II34901);
  not NOT_10634(II34909,g26265);
  not NOT_10635(g26788,II34909);
  not NOT_10636(II34916,g26240);
  not NOT_10637(g26793,II34916);
  not NOT_10638(II34921,g26217);
  not NOT_10639(g26796,II34921);
  not NOT_10640(II34946,g26534);
  not NOT_10641(g26819,II34946);
  not NOT_10642(II34957,g26541);
  not NOT_10643(g26828,II34957);
  not NOT_10644(II34961,g26545);
  not NOT_10645(g26830,II34961);
  not NOT_10646(II34964,g26547);
  not NOT_10647(g26831,II34964);
  not NOT_10648(II34967,g26553);
  not NOT_10649(g26832,II34967);
  not NOT_10650(II34971,g26557);
  not NOT_10651(g26834,II34971);
  not NOT_10652(II34974,g26168);
  not NOT_10653(g26835,II34974);
  not NOT_10654(II34977,g26559);
  not NOT_10655(g26836,II34977);
  not NOT_10656(II34980,g26458);
  not NOT_10657(g26837,II34980);
  not NOT_10658(II34983,g26569);
  not NOT_10659(g26840,II34983);
  not NOT_10660(II34986,g26160);
  not NOT_10661(g26841,II34986);
  not NOT_10662(II34990,g26573);
  not NOT_10663(g26843,II34990);
  not NOT_10664(II34993,g26575);
  not NOT_10665(g26844,II34993);
  not NOT_10666(II34997,g26482);
  not NOT_10667(g26846,II34997);
  not NOT_10668(II35000,g26336);
  not NOT_10669(g26849,II35000);
  not NOT_10670(II35003,g26592);
  not NOT_10671(g26850,II35003);
  not NOT_10672(II35007,g26596);
  not NOT_10673(g26852,II35007);
  not NOT_10674(II35011,g26304);
  not NOT_10675(g26854,II35011);
  not NOT_10676(II35014,g26498);
  not NOT_10677(g26855,II35014);
  not NOT_10678(II35017,g26616);
  not NOT_10679(g26858,II35017);
  not NOT_10680(II35028,g26513);
  not NOT_10681(g26861,II35028);
  not NOT_10682(II35031,g26529);
  not NOT_10683(g26864,II35031);
  not NOT_10684(II35049,g26530);
  not NOT_10685(g26868,II35049);
  not NOT_10686(II35053,g26655);
  not NOT_10687(g26872,II35053);
  not NOT_10688(II35064,g26531);
  not NOT_10689(g26875,II35064);
  not NOT_10690(II35067,g26659);
  not NOT_10691(g26876,II35067);
  not NOT_10692(II35072,g26661);
  not NOT_10693(g26881,II35072);
  not NOT_10694(II35076,g26532);
  not NOT_10695(g26883,II35076);
  not NOT_10696(II35079,g26664);
  not NOT_10697(g26884,II35079);
  not NOT_10698(II35083,g26665);
  not NOT_10699(g26886,II35083);
  not NOT_10700(II35087,g26667);
  not NOT_10701(g26890,II35087);
  not NOT_10702(II35092,g26669);
  not NOT_10703(g26895,II35092);
  not NOT_10704(II35095,g26670);
  not NOT_10705(g26896,II35095);
  not NOT_10706(II35099,g26672);
  not NOT_10707(g26900,II35099);
  not NOT_10708(II35106,g26675);
  not NOT_10709(g26909,II35106);
  not NOT_10710(II35109,g26676);
  not NOT_10711(g26910,II35109);
  not NOT_10712(II35116,g26025);
  not NOT_10713(g26921,II35116);
  not NOT_10714(g26922,g26283);
  not NOT_10715(g26935,g26327);
  not NOT_10716(g26944,g26374);
  not NOT_10717(g26950,g26417);
  not NOT_10718(II35136,g26660);
  not NOT_10719(g26953,II35136);
  not NOT_10720(g26954,g26549);
  not NOT_10721(II35141,g26666);
  not NOT_10722(g26956,II35141);
  not NOT_10723(g26957,g26577);
  not NOT_10724(II35146,g26671);
  not NOT_10725(g26959,II35146);
  not NOT_10726(g26960,g26597);
  not NOT_10727(II35153,g26677);
  not NOT_10728(g26964,II35153);
  not NOT_10729(II35172,g26272);
  not NOT_10730(g26983,II35172);
  not NOT_10731(g26987,g26056);
  not NOT_10732(g27010,g26063);
  not NOT_10733(g27036,g26070);
  not NOT_10734(g27064,g26076);
  not NOT_10735(II35254,g26048);
  not NOT_10736(g27075,II35254);
  not NOT_10737(II35283,g26031);
  not NOT_10738(g27102,II35283);
  not NOT_10739(II35297,g26199);
  not NOT_10740(g27114,II35297);
  not NOT_10741(II35301,g26037);
  not NOT_10742(g27116,II35301);
  not NOT_10743(II35313,g26534);
  not NOT_10744(g27126,II35313);
  not NOT_10745(II35319,g26183);
  not NOT_10746(g27132,II35319);
  not NOT_10747(g27133,g26105);
  not NOT_10748(g27134,g26175);
  not NOT_10749(g27135,g26178);
  not NOT_10750(g27136,g26196);
  not NOT_10751(g27137,g26202);
  not NOT_10752(g27138,g26223);
  not NOT_10753(g27139,g26226);
  not NOT_10754(g27140,g26136);
  not NOT_10755(g27141,g26251);
  not NOT_10756(g27142,g26254);
  not NOT_10757(g27143,g26150);
  not NOT_10758(II35334,g26106);
  not NOT_10759(g27145,II35334);
  not NOT_10760(g27146,g26358);
  not NOT_10761(g27148,g26393);
  not NOT_10762(II35341,g26120);
  not NOT_10763(g27150,II35341);
  not NOT_10764(g27151,g26401);
  not NOT_10765(g27153,g26429);
  not NOT_10766(II35347,g26265);
  not NOT_10767(g27154,II35347);
  not NOT_10768(g27155,g26434);
  not NOT_10769(II35351,g26272);
  not NOT_10770(g27156,II35351);
  not NOT_10771(II35355,g26130);
  not NOT_10772(g27158,II35355);
  not NOT_10773(g27159,g26442);
  not NOT_10774(II35360,g26295);
  not NOT_10775(g27161,II35360);
  not NOT_10776(g27162,g26461);
  not NOT_10777(II35364,g26304);
  not NOT_10778(g27163,II35364);
  not NOT_10779(g27164,g26466);
  not NOT_10780(II35369,g26144);
  not NOT_10781(g27166,II35369);
  not NOT_10782(g27167,g26474);
  not NOT_10783(II35373,g26189);
  not NOT_10784(g27168,II35373);
  not NOT_10785(II35376,g26336);
  not NOT_10786(g27171,II35376);
  not NOT_10787(g27172,g26485);
  not NOT_10788(g27173,g26490);
  not NOT_10789(II35383,g26160);
  not NOT_10790(g27176,II35383);
  not NOT_10791(g27177,g26501);
  not NOT_10792(II35389,g26168);
  not NOT_10793(g27180,II35389);
  not NOT_10794(II35394,g26183);
  not NOT_10795(g27183,II35394);
  not NOT_10796(II35399,g26199);
  not NOT_10797(g27186,II35399);
  not NOT_10798(II35404,g26864);
  not NOT_10799(g27189,II35404);
  not NOT_10800(II35407,g27145);
  not NOT_10801(g27190,II35407);
  not NOT_10802(II35410,g26872);
  not NOT_10803(g27191,II35410);
  not NOT_10804(II35413,g26876);
  not NOT_10805(g27192,II35413);
  not NOT_10806(II35416,g26884);
  not NOT_10807(g27193,II35416);
  not NOT_10808(II35419,g26828);
  not NOT_10809(g27194,II35419);
  not NOT_10810(II35422,g26830);
  not NOT_10811(g27195,II35422);
  not NOT_10812(II35425,g26832);
  not NOT_10813(g27196,II35425);
  not NOT_10814(II35428,g26953);
  not NOT_10815(g27197,II35428);
  not NOT_10816(II35431,g26868);
  not NOT_10817(g27198,II35431);
  not NOT_10818(II35434,g27150);
  not NOT_10819(g27199,II35434);
  not NOT_10820(II35437,g27183);
  not NOT_10821(g27200,II35437);
  not NOT_10822(II35440,g27186);
  not NOT_10823(g27201,II35440);
  not NOT_10824(II35443,g26757);
  not NOT_10825(g27202,II35443);
  not NOT_10826(II35446,g26762);
  not NOT_10827(g27203,II35446);
  not NOT_10828(II35449,g27154);
  not NOT_10829(g27204,II35449);
  not NOT_10830(II35452,g27161);
  not NOT_10831(g27205,II35452);
  not NOT_10832(II35455,g26881);
  not NOT_10833(g27206,II35455);
  not NOT_10834(II35458,g26886);
  not NOT_10835(g27207,II35458);
  not NOT_10836(II35461,g26895);
  not NOT_10837(g27208,II35461);
  not NOT_10838(II35464,g26831);
  not NOT_10839(g27209,II35464);
  not NOT_10840(II35467,g26834);
  not NOT_10841(g27210,II35467);
  not NOT_10842(II35470,g26840);
  not NOT_10843(g27211,II35470);
  not NOT_10844(II35473,g27156);
  not NOT_10845(g27212,II35473);
  not NOT_10846(II35476,g27163);
  not NOT_10847(g27213,II35476);
  not NOT_10848(II35479,g27171);
  not NOT_10849(g27214,II35479);
  not NOT_10850(II35482,g27176);
  not NOT_10851(g27215,II35482);
  not NOT_10852(II35485,g27180);
  not NOT_10853(g27216,II35485);
  not NOT_10854(II35488,g26819);
  not NOT_10855(g27217,II35488);
  not NOT_10856(II35491,g26956);
  not NOT_10857(g27218,II35491);
  not NOT_10858(II35494,g26875);
  not NOT_10859(g27219,II35494);
  not NOT_10860(II35497,g27158);
  not NOT_10861(g27220,II35497);
  not NOT_10862(II35500,g26890);
  not NOT_10863(g27221,II35500);
  not NOT_10864(II35503,g26896);
  not NOT_10865(g27222,II35503);
  not NOT_10866(II35506,g26909);
  not NOT_10867(g27223,II35506);
  not NOT_10868(II35509,g26836);
  not NOT_10869(g27224,II35509);
  not NOT_10870(II35512,g26843);
  not NOT_10871(g27225,II35512);
  not NOT_10872(II35515,g26850);
  not NOT_10873(g27226,II35515);
  not NOT_10874(II35518,g26959);
  not NOT_10875(g27227,II35518);
  not NOT_10876(II35521,g26883);
  not NOT_10877(g27228,II35521);
  not NOT_10878(II35524,g27166);
  not NOT_10879(g27229,II35524);
  not NOT_10880(II35527,g26900);
  not NOT_10881(g27230,II35527);
  not NOT_10882(II35530,g26910);
  not NOT_10883(g27231,II35530);
  not NOT_10884(II35533,g26921);
  not NOT_10885(g27232,II35533);
  not NOT_10886(II35536,g26844);
  not NOT_10887(g27233,II35536);
  not NOT_10888(II35539,g26852);
  not NOT_10889(g27234,II35539);
  not NOT_10890(II35542,g26858);
  not NOT_10891(g27235,II35542);
  not NOT_10892(II35545,g26964);
  not NOT_10893(g27236,II35545);
  not NOT_10894(II35548,g27116);
  not NOT_10895(g27237,II35548);
  not NOT_10896(II35551,g27075);
  not NOT_10897(g27238,II35551);
  not NOT_10898(II35554,g27102);
  not NOT_10899(g27239,II35554);
  not NOT_10900(g27349,g27126);
  not NOT_10901(II35667,g27120);
  not NOT_10902(g27353,II35667);
  not NOT_10903(II35673,g27123);
  not NOT_10904(g27357,II35673);
  not NOT_10905(II35678,g27129);
  not NOT_10906(g27360,II35678);
  not NOT_10907(II35681,g26869);
  not NOT_10908(g27361,II35681);
  not NOT_10909(II35686,g27131);
  not NOT_10910(g27366,II35686);
  not NOT_10911(II35689,g26878);
  not NOT_10912(g27367,II35689);
  not NOT_10913(II35695,g26887);
  not NOT_10914(g27373,II35695);
  not NOT_10915(II35698,g26897);
  not NOT_10916(g27376,II35698);
  not NOT_10917(II35708,g26974);
  not NOT_10918(g27380,II35708);
  not NOT_10919(II35711,g26974);
  not NOT_10920(g27381,II35711);
  not NOT_10921(g27383,g27133);
  not NOT_10922(g27384,g27140);
  not NOT_10923(II35723,g27168);
  not NOT_10924(g27385,II35723);
  not NOT_10925(g27386,g27143);
  not NOT_10926(II35727,g26902);
  not NOT_10927(g27387,II35727);
  not NOT_10928(II35731,g26892);
  not NOT_10929(g27391,II35731);
  not NOT_10930(II35737,g26915);
  not NOT_10931(g27397,II35737);
  not NOT_10932(II35741,g27118);
  not NOT_10933(g27401,II35741);
  not NOT_10934(II35744,g26906);
  not NOT_10935(g27404,II35744);
  not NOT_10936(II35750,g26928);
  not NOT_10937(g27410,II35750);
  not NOT_10938(II35756,g27117);
  not NOT_10939(g27416,II35756);
  not NOT_10940(II35759,g27121);
  not NOT_10941(g27419,II35759);
  not NOT_10942(II35762,g26918);
  not NOT_10943(g27422,II35762);
  not NOT_10944(II35768,g26941);
  not NOT_10945(g27428,II35768);
  not NOT_10946(II35772,g26772);
  not NOT_10947(g27432,II35772);
  not NOT_10948(II35777,g27119);
  not NOT_10949(g27437,II35777);
  not NOT_10950(II35780,g27124);
  not NOT_10951(g27440,II35780);
  not NOT_10952(II35783,g26931);
  not NOT_10953(g27443,II35783);
  not NOT_10954(g27449,g26837);
  not NOT_10955(II35791,g26779);
  not NOT_10956(g27451,II35791);
  not NOT_10957(II35796,g27122);
  not NOT_10958(g27456,II35796);
  not NOT_10959(II35799,g27130);
  not NOT_10960(g27459,II35799);
  not NOT_10961(II35803,g26803);
  not NOT_10962(g27463,II35803);
  not NOT_10963(g27465,g26846);
  not NOT_10964(II35809,g26785);
  not NOT_10965(g27467,II35809);
  not NOT_10966(II35814,g27125);
  not NOT_10967(g27472,II35814);
  not NOT_10968(II35817,g26922);
  not NOT_10969(g27475,II35817);
  not NOT_10970(II35821,g26804);
  not NOT_10971(g27479,II35821);
  not NOT_10972(II35824,g26805);
  not NOT_10973(g27480,II35824);
  not NOT_10974(II35829,g26806);
  not NOT_10975(g27483,II35829);
  not NOT_10976(g27484,g26855);
  not NOT_10977(II35834,g26792);
  not NOT_10978(g27486,II35834);
  not NOT_10979(II35837,g26911);
  not NOT_10980(g27489,II35837);
  not NOT_10981(II35841,g26807);
  not NOT_10982(g27493,II35841);
  not NOT_10983(II35844,g26808);
  not NOT_10984(g27494,II35844);
  not NOT_10985(II35849,g26776);
  not NOT_10986(g27497,II35849);
  not NOT_10987(II35852,g26935);
  not NOT_10988(g27498,II35852);
  not NOT_10989(II35856,g26809);
  not NOT_10990(g27502,II35856);
  not NOT_10991(II35859,g26810);
  not NOT_10992(g27503,II35859);
  not NOT_10993(II35863,g26811);
  not NOT_10994(g27505,II35863);
  not NOT_10995(g27506,g26861);
  not NOT_10996(II35868,g26812);
  not NOT_10997(g27508,II35868);
  not NOT_10998(II35872,g26925);
  not NOT_10999(g27510,II35872);
  not NOT_11000(II35876,g26813);
  not NOT_11001(g27514,II35876);
  not NOT_11002(II35879,g26814);
  not NOT_11003(g27515,II35879);
  not NOT_11004(II35883,g26781);
  not NOT_11005(g27517,II35883);
  not NOT_11006(II35886,g26944);
  not NOT_11007(g27518,II35886);
  not NOT_11008(II35890,g26815);
  not NOT_11009(g27522,II35890);
  not NOT_11010(II35893,g26816);
  not NOT_11011(g27523,II35893);
  not NOT_11012(II35897,g26817);
  not NOT_11013(g27525,II35897);
  not NOT_11014(II35900,g26786);
  not NOT_11015(g27526,II35900);
  not NOT_11016(II35915,g26818);
  not NOT_11017(g27533,II35915);
  not NOT_11018(II35919,g26938);
  not NOT_11019(g27535,II35919);
  not NOT_11020(II35923,g26820);
  not NOT_11021(g27539,II35923);
  not NOT_11022(II35926,g26821);
  not NOT_11023(g27540,II35926);
  not NOT_11024(II35930,g26789);
  not NOT_11025(g27542,II35930);
  not NOT_11026(II35933,g26950);
  not NOT_11027(g27543,II35933);
  not NOT_11028(II35937,g26822);
  not NOT_11029(g27547,II35937);
  not NOT_11030(II35940,g26823);
  not NOT_11031(g27548,II35940);
  not NOT_11032(II35953,g26824);
  not NOT_11033(g27553,II35953);
  not NOT_11034(II35957,g26947);
  not NOT_11035(g27555,II35957);
  not NOT_11036(II35961,g26825);
  not NOT_11037(g27559,II35961);
  not NOT_11038(II35964,g26826);
  not NOT_11039(g27560,II35964);
  not NOT_11040(II35968,g26795);
  not NOT_11041(g27562,II35968);
  not NOT_11042(II35983,g26827);
  not NOT_11043(g27569,II35983);
  not NOT_11044(II36008,g26798);
  not NOT_11045(g27586,II36008);
  not NOT_11046(g27589,g27168);
  not NOT_11047(g27590,g27144);
  not NOT_11048(g27595,g27149);
  not NOT_11049(g27599,g27147);
  not NOT_11050(g27604,g27157);
  not NOT_11051(g27608,g27152);
  not NOT_11052(g27613,g27165);
  not NOT_11053(g27617,g27160);
  not NOT_11054(g27622,g27174);
  not NOT_11055(II36032,g27113);
  not NOT_11056(g27632,II36032);
  not NOT_11057(II36042,g26960);
  not NOT_11058(g27662,II36042);
  not NOT_11059(II36046,g26957);
  not NOT_11060(g27667,II36046);
  not NOT_11061(II36052,g26954);
  not NOT_11062(g27674,II36052);
  not NOT_11063(II36060,g27353);
  not NOT_11064(g27683,II36060);
  not NOT_11065(II36063,g27463);
  not NOT_11066(g27684,II36063);
  not NOT_11067(II36066,g27479);
  not NOT_11068(g27685,II36066);
  not NOT_11069(II36069,g27493);
  not NOT_11070(g27686,II36069);
  not NOT_11071(II36072,g27480);
  not NOT_11072(g27687,II36072);
  not NOT_11073(II36075,g27494);
  not NOT_11074(g27688,II36075);
  not NOT_11075(II36078,g27508);
  not NOT_11076(g27689,II36078);
  not NOT_11077(II36081,g27497);
  not NOT_11078(g27690,II36081);
  not NOT_11079(II36084,g27357);
  not NOT_11080(g27691,II36084);
  not NOT_11081(II36087,g27483);
  not NOT_11082(g27692,II36087);
  not NOT_11083(II36090,g27502);
  not NOT_11084(g27693,II36090);
  not NOT_11085(II36093,g27514);
  not NOT_11086(g27694,II36093);
  not NOT_11087(II36096,g27503);
  not NOT_11088(g27695,II36096);
  not NOT_11089(II36099,g27515);
  not NOT_11090(g27696,II36099);
  not NOT_11091(II36102,g27533);
  not NOT_11092(g27697,II36102);
  not NOT_11093(II36105,g27517);
  not NOT_11094(g27698,II36105);
  not NOT_11095(II36108,g27360);
  not NOT_11096(g27699,II36108);
  not NOT_11097(II36111,g27505);
  not NOT_11098(g27700,II36111);
  not NOT_11099(II36114,g27522);
  not NOT_11100(g27701,II36114);
  not NOT_11101(II36117,g27539);
  not NOT_11102(g27702,II36117);
  not NOT_11103(II36120,g27523);
  not NOT_11104(g27703,II36120);
  not NOT_11105(II36123,g27540);
  not NOT_11106(g27704,II36123);
  not NOT_11107(II36126,g27553);
  not NOT_11108(g27705,II36126);
  not NOT_11109(II36129,g27542);
  not NOT_11110(g27706,II36129);
  not NOT_11111(II36132,g27366);
  not NOT_11112(g27707,II36132);
  not NOT_11113(II36135,g27525);
  not NOT_11114(g27708,II36135);
  not NOT_11115(II36138,g27547);
  not NOT_11116(g27709,II36138);
  not NOT_11117(II36141,g27559);
  not NOT_11118(g27710,II36141);
  not NOT_11119(II36144,g27548);
  not NOT_11120(g27711,II36144);
  not NOT_11121(II36147,g27560);
  not NOT_11122(g27712,II36147);
  not NOT_11123(II36150,g27569);
  not NOT_11124(g27713,II36150);
  not NOT_11125(II36153,g27562);
  not NOT_11126(g27714,II36153);
  not NOT_11127(II36156,g27586);
  not NOT_11128(g27715,II36156);
  not NOT_11129(II36159,g27526);
  not NOT_11130(g27716,II36159);
  not NOT_11131(II36162,g27385);
  not NOT_11132(g27717,II36162);
  not NOT_11133(g27748,g27632);
  not NOT_11134(II36213,g27571);
  not NOT_11135(g27776,II36213);
  not NOT_11136(II36217,g27580);
  not NOT_11137(g27780,II36217);
  not NOT_11138(II36221,g27662);
  not NOT_11139(g27784,II36221);
  not NOT_11140(II36224,g27589);
  not NOT_11141(g27785,II36224);
  not NOT_11142(II36227,g27594);
  not NOT_11143(g27786,II36227);
  not NOT_11144(II36230,g27583);
  not NOT_11145(g27787,II36230);
  not NOT_11146(II36234,g27667);
  not NOT_11147(g27791,II36234);
  not NOT_11148(II36237,g27662);
  not NOT_11149(g27792,II36237);
  not NOT_11150(II36240,g27603);
  not NOT_11151(g27793,II36240);
  not NOT_11152(II36243,g27587);
  not NOT_11153(g27794,II36243);
  not NOT_11154(II36246,g27674);
  not NOT_11155(g27797,II36246);
  not NOT_11156(II36250,g27612);
  not NOT_11157(g27799,II36250);
  not NOT_11158(II36253,g27674);
  not NOT_11159(g27800,II36253);
  not NOT_11160(II36264,g27621);
  not NOT_11161(g27805,II36264);
  not NOT_11162(II36267,g27395);
  not NOT_11163(g27806,II36267);
  not NOT_11164(II36280,g27390);
  not NOT_11165(g27817,II36280);
  not NOT_11166(II36283,g27408);
  not NOT_11167(g27820,II36283);
  not NOT_11168(II36296,g27626);
  not NOT_11169(g27831,II36296);
  not NOT_11170(II36307,g27400);
  not NOT_11171(g27839,II36307);
  not NOT_11172(II36311,g27426);
  not NOT_11173(g27843,II36311);
  not NOT_11174(II36321,g27627);
  not NOT_11175(g27847,II36321);
  not NOT_11176(II36327,g27413);
  not NOT_11177(g27858,II36327);
  not NOT_11178(II36330,g27447);
  not NOT_11179(g27861,II36330);
  not NOT_11180(II36337,g27628);
  not NOT_11181(g27872,II36337);
  not NOT_11182(II36341,g27431);
  not NOT_11183(g27879,II36341);
  not NOT_11184(II36347,g27630);
  not NOT_11185(g27889,II36347);
  not NOT_11186(II36354,g27662);
  not NOT_11187(g27903,II36354);
  not NOT_11188(II36358,g27672);
  not NOT_11189(g27905,II36358);
  not NOT_11190(II36362,g27667);
  not NOT_11191(g27907,II36362);
  not NOT_11192(II36367,g27678);
  not NOT_11193(g27910,II36367);
  not NOT_11194(II36371,g27674);
  not NOT_11195(g27912,II36371);
  not NOT_11196(II36379,g27682);
  not NOT_11197(g27918,II36379);
  not NOT_11198(II36382,g27563);
  not NOT_11199(g27919,II36382);
  not NOT_11200(II36390,g27243);
  not NOT_11201(g27927,II36390);
  not NOT_11202(II36393,g27572);
  not NOT_11203(g27928,II36393);
  not NOT_11204(II36397,g27574);
  not NOT_11205(g27932,II36397);
  not NOT_11206(II36404,g27450);
  not NOT_11207(g27939,II36404);
  not NOT_11208(II36407,g27581);
  not NOT_11209(g27942,II36407);
  not NOT_11210(II36411,g27582);
  not NOT_11211(g27946,II36411);
  not NOT_11212(II36417,g27462);
  not NOT_11213(g27952,II36417);
  not NOT_11214(II36420,g27253);
  not NOT_11215(g27955,II36420);
  not NOT_11216(II36423,g27466);
  not NOT_11217(g27956,II36423);
  not NOT_11218(II36426,g27584);
  not NOT_11219(g27959,II36426);
  not NOT_11220(II36432,g27585);
  not NOT_11221(g27965,II36432);
  not NOT_11222(g27969,g27361);
  not NOT_11223(II36438,g27255);
  not NOT_11224(g27971,II36438);
  not NOT_11225(II36441,g27256);
  not NOT_11226(g27972,II36441);
  not NOT_11227(II36444,g27482);
  not NOT_11228(g27973,II36444);
  not NOT_11229(II36447,g27257);
  not NOT_11230(g27976,II36447);
  not NOT_11231(II36450,g27485);
  not NOT_11232(g27977,II36450);
  not NOT_11233(II36454,g27588);
  not NOT_11234(g27981,II36454);
  not NOT_11235(II36459,g27258);
  not NOT_11236(g27986,II36459);
  not NOT_11237(II36462,g27259);
  not NOT_11238(g27987,II36462);
  not NOT_11239(II36465,g27260);
  not NOT_11240(g27988,II36465);
  not NOT_11241(II36468,g27261);
  not NOT_11242(g27989,II36468);
  not NOT_11243(g27990,g27367);
  not NOT_11244(II36473,g27262);
  not NOT_11245(g27992,II36473);
  not NOT_11246(II36476,g27263);
  not NOT_11247(g27993,II36476);
  not NOT_11248(II36479,g27504);
  not NOT_11249(g27994,II36479);
  not NOT_11250(II36483,g27264);
  not NOT_11251(g27998,II36483);
  not NOT_11252(II36486,g27507);
  not NOT_11253(g27999,II36486);
  not NOT_11254(II36490,g27265);
  not NOT_11255(g28003,II36490);
  not NOT_11256(II36493,g27266);
  not NOT_11257(g28004,II36493);
  not NOT_11258(II36496,g27267);
  not NOT_11259(g28005,II36496);
  not NOT_11260(II36499,g27268);
  not NOT_11261(g28006,II36499);
  not NOT_11262(II36502,g27269);
  not NOT_11263(g28007,II36502);
  not NOT_11264(II36507,g27270);
  not NOT_11265(g28010,II36507);
  not NOT_11266(II36510,g27271);
  not NOT_11267(g28011,II36510);
  not NOT_11268(II36513,g27272);
  not NOT_11269(g28012,II36513);
  not NOT_11270(II36516,g27273);
  not NOT_11271(g28013,II36516);
  not NOT_11272(g28014,g27373);
  not NOT_11273(II36521,g27274);
  not NOT_11274(g28016,II36521);
  not NOT_11275(II36524,g27275);
  not NOT_11276(g28017,II36524);
  not NOT_11277(II36527,g27524);
  not NOT_11278(g28018,II36527);
  not NOT_11279(II36530,g27276);
  not NOT_11280(g28021,II36530);
  not NOT_11281(II36533,g27277);
  not NOT_11282(g28022,II36533);
  not NOT_11283(II36536,g27278);
  not NOT_11284(g28023,II36536);
  not NOT_11285(II36539,g27279);
  not NOT_11286(g28024,II36539);
  not NOT_11287(II36542,g27280);
  not NOT_11288(g28025,II36542);
  not NOT_11289(II36545,g27281);
  not NOT_11290(g28026,II36545);
  not NOT_11291(II36551,g27282);
  not NOT_11292(g28030,II36551);
  not NOT_11293(II36554,g27283);
  not NOT_11294(g28031,II36554);
  not NOT_11295(II36557,g27284);
  not NOT_11296(g28032,II36557);
  not NOT_11297(II36560,g27285);
  not NOT_11298(g28033,II36560);
  not NOT_11299(II36563,g27286);
  not NOT_11300(g28034,II36563);
  not NOT_11301(II36568,g27287);
  not NOT_11302(g28037,II36568);
  not NOT_11303(II36571,g27288);
  not NOT_11304(g28038,II36571);
  not NOT_11305(II36574,g27289);
  not NOT_11306(g28039,II36574);
  not NOT_11307(II36577,g27290);
  not NOT_11308(g28040,II36577);
  not NOT_11309(g28041,g27376);
  not NOT_11310(II36582,g27291);
  not NOT_11311(g28043,II36582);
  not NOT_11312(II36585,g27292);
  not NOT_11313(g28044,II36585);
  not NOT_11314(II36588,g27293);
  not NOT_11315(g28045,II36588);
  not NOT_11316(II36598,g27294);
  not NOT_11317(g28047,II36598);
  not NOT_11318(II36601,g27295);
  not NOT_11319(g28048,II36601);
  not NOT_11320(II36604,g27296);
  not NOT_11321(g28049,II36604);
  not NOT_11322(II36609,g27297);
  not NOT_11323(g28052,II36609);
  not NOT_11324(II36612,g27298);
  not NOT_11325(g28053,II36612);
  not NOT_11326(II36615,g27299);
  not NOT_11327(g28054,II36615);
  not NOT_11328(II36618,g27300);
  not NOT_11329(g28055,II36618);
  not NOT_11330(II36621,g27301);
  not NOT_11331(g28056,II36621);
  not NOT_11332(II36627,g27302);
  not NOT_11333(g28060,II36627);
  not NOT_11334(II36630,g27303);
  not NOT_11335(g28061,II36630);
  not NOT_11336(II36633,g27304);
  not NOT_11337(g28062,II36633);
  not NOT_11338(II36636,g27305);
  not NOT_11339(g28063,II36636);
  not NOT_11340(II36639,g27306);
  not NOT_11341(g28064,II36639);
  not NOT_11342(II36644,g27307);
  not NOT_11343(g28067,II36644);
  not NOT_11344(II36647,g27308);
  not NOT_11345(g28068,II36647);
  not NOT_11346(II36650,g27309);
  not NOT_11347(g28069,II36650);
  not NOT_11348(II36653,g27310);
  not NOT_11349(g28070,II36653);
  not NOT_11350(II36656,g27311);
  not NOT_11351(g28071,II36656);
  not NOT_11352(II36659,g27312);
  not NOT_11353(g28072,II36659);
  not NOT_11354(II36663,g27313);
  not NOT_11355(g28074,II36663);
  not NOT_11356(II36673,g27314);
  not NOT_11357(g28076,II36673);
  not NOT_11358(II36676,g27315);
  not NOT_11359(g28077,II36676);
  not NOT_11360(II36679,g27316);
  not NOT_11361(g28078,II36679);
  not NOT_11362(II36684,g27317);
  not NOT_11363(g28081,II36684);
  not NOT_11364(II36687,g27318);
  not NOT_11365(g28082,II36687);
  not NOT_11366(II36690,g27319);
  not NOT_11367(g28083,II36690);
  not NOT_11368(II36693,g27320);
  not NOT_11369(g28084,II36693);
  not NOT_11370(II36696,g27321);
  not NOT_11371(g28085,II36696);
  not NOT_11372(II36702,g27322);
  not NOT_11373(g28089,II36702);
  not NOT_11374(II36705,g27323);
  not NOT_11375(g28090,II36705);
  not NOT_11376(II36708,g27324);
  not NOT_11377(g28091,II36708);
  not NOT_11378(II36711,g27325);
  not NOT_11379(g28092,II36711);
  not NOT_11380(II36714,g27326);
  not NOT_11381(g28093,II36714);
  not NOT_11382(II36718,g27327);
  not NOT_11383(g28095,II36718);
  not NOT_11384(II36721,g27328);
  not NOT_11385(g28096,II36721);
  not NOT_11386(II36724,g27329);
  not NOT_11387(g28097,II36724);
  not NOT_11388(II36728,g27330);
  not NOT_11389(g28099,II36728);
  not NOT_11390(II36738,g27331);
  not NOT_11391(g28101,II36738);
  not NOT_11392(II36741,g27332);
  not NOT_11393(g28102,II36741);
  not NOT_11394(II36744,g27333);
  not NOT_11395(g28103,II36744);
  not NOT_11396(II36749,g27334);
  not NOT_11397(g28106,II36749);
  not NOT_11398(II36752,g27335);
  not NOT_11399(g28107,II36752);
  not NOT_11400(II36755,g27336);
  not NOT_11401(g28108,II36755);
  not NOT_11402(II36758,g27337);
  not NOT_11403(g28109,II36758);
  not NOT_11404(II36761,g27338);
  not NOT_11405(g28110,II36761);
  not NOT_11406(II36766,g27339);
  not NOT_11407(g28113,II36766);
  not NOT_11408(II36769,g27340);
  not NOT_11409(g28114,II36769);
  not NOT_11410(II36772,g27341);
  not NOT_11411(g28115,II36772);
  not NOT_11412(II36776,g27342);
  not NOT_11413(g28117,II36776);
  not NOT_11414(II36786,g27343);
  not NOT_11415(g28119,II36786);
  not NOT_11416(II36789,g27344);
  not NOT_11417(g28120,II36789);
  not NOT_11418(II36792,g27345);
  not NOT_11419(g28121,II36792);
  not NOT_11420(II36797,g27346);
  not NOT_11421(g28124,II36797);
  not NOT_11422(II36800,g27347);
  not NOT_11423(g28125,II36800);
  not NOT_11424(II36803,g27348);
  not NOT_11425(g28126,II36803);
  not NOT_11426(g28128,g27528);
  not NOT_11427(II36808,g27354);
  not NOT_11428(g28132,II36808);
  not NOT_11429(g28133,g27550);
  not NOT_11430(g28137,g27566);
  not NOT_11431(g28141,g27576);
  not NOT_11432(g28149,g27667);
  not NOT_11433(g28150,g27387);
  not NOT_11434(g28151,g27381);
  not NOT_11435(g28152,g27391);
  not NOT_11436(g28153,g27397);
  not NOT_11437(g28154,g27401);
  not NOT_11438(g28155,g27404);
  not NOT_11439(g28156,g27410);
  not NOT_11440(g28158,g27416);
  not NOT_11441(g28159,g27419);
  not NOT_11442(g28160,g27422);
  not NOT_11443(g28161,g27428);
  not NOT_11444(g28162,g27432);
  not NOT_11445(g28163,g27437);
  not NOT_11446(g28164,g27440);
  not NOT_11447(g28165,g27443);
  not NOT_11448(g28166,g27451);
  not NOT_11449(g28167,g27456);
  not NOT_11450(g28168,g27459);
  not NOT_11451(g28169,g27467);
  not NOT_11452(g28170,g27472);
  not NOT_11453(g28172,g27475);
  not NOT_11454(g28173,g27486);
  not NOT_11455(g28174,g27489);
  not NOT_11456(g28175,g27498);
  not NOT_11457(g28177,g27510);
  not NOT_11458(g28178,g27518);
  not NOT_11459(II36848,g27383);
  not NOT_11460(g28179,II36848);
  not NOT_11461(g28186,g27535);
  not NOT_11462(g28187,g27543);
  not NOT_11463(g28190,g27555);
  not NOT_11464(II36860,g27386);
  not NOT_11465(g28194,II36860);
  not NOT_11466(II36864,g27384);
  not NOT_11467(g28200,II36864);
  not NOT_11468(II36867,g27786);
  not NOT_11469(g28206,II36867);
  not NOT_11470(II36870,g27955);
  not NOT_11471(g28207,II36870);
  not NOT_11472(II36873,g27971);
  not NOT_11473(g28208,II36873);
  not NOT_11474(II36876,g27986);
  not NOT_11475(g28209,II36876);
  not NOT_11476(II36879,g27972);
  not NOT_11477(g28210,II36879);
  not NOT_11478(II36882,g27987);
  not NOT_11479(g28211,II36882);
  not NOT_11480(II36885,g28003);
  not NOT_11481(g28212,II36885);
  not NOT_11482(II36888,g27988);
  not NOT_11483(g28213,II36888);
  not NOT_11484(II36891,g28004);
  not NOT_11485(g28214,II36891);
  not NOT_11486(II36894,g28022);
  not NOT_11487(g28215,II36894);
  not NOT_11488(II36897,g28005);
  not NOT_11489(g28216,II36897);
  not NOT_11490(II36900,g28023);
  not NOT_11491(g28217,II36900);
  not NOT_11492(II36903,g28045);
  not NOT_11493(g28218,II36903);
  not NOT_11494(II36906,g27989);
  not NOT_11495(g28219,II36906);
  not NOT_11496(II36909,g28006);
  not NOT_11497(g28220,II36909);
  not NOT_11498(II36912,g28024);
  not NOT_11499(g28221,II36912);
  not NOT_11500(II36915,g28007);
  not NOT_11501(g28222,II36915);
  not NOT_11502(II36918,g28025);
  not NOT_11503(g28223,II36918);
  not NOT_11504(II36921,g28047);
  not NOT_11505(g28224,II36921);
  not NOT_11506(II36924,g28026);
  not NOT_11507(g28225,II36924);
  not NOT_11508(II36927,g28048);
  not NOT_11509(g28226,II36927);
  not NOT_11510(II36930,g28071);
  not NOT_11511(g28227,II36930);
  not NOT_11512(II36933,g28049);
  not NOT_11513(g28228,II36933);
  not NOT_11514(II36936,g28072);
  not NOT_11515(g28229,II36936);
  not NOT_11516(II36939,g28095);
  not NOT_11517(g28230,II36939);
  not NOT_11518(II36942,g27905);
  not NOT_11519(g28231,II36942);
  not NOT_11520(II36945,g27793);
  not NOT_11521(g28232,II36945);
  not NOT_11522(II36948,g27976);
  not NOT_11523(g28233,II36948);
  not NOT_11524(II36951,g27992);
  not NOT_11525(g28234,II36951);
  not NOT_11526(II36954,g28010);
  not NOT_11527(g28235,II36954);
  not NOT_11528(II36957,g27993);
  not NOT_11529(g28236,II36957);
  not NOT_11530(II36960,g28011);
  not NOT_11531(g28237,II36960);
  not NOT_11532(II36963,g28030);
  not NOT_11533(g28238,II36963);
  not NOT_11534(II36966,g28012);
  not NOT_11535(g28239,II36966);
  not NOT_11536(II36969,g28031);
  not NOT_11537(g28240,II36969);
  not NOT_11538(II36972,g28052);
  not NOT_11539(g28241,II36972);
  not NOT_11540(II36975,g28032);
  not NOT_11541(g28242,II36975);
  not NOT_11542(II36978,g28053);
  not NOT_11543(g28243,II36978);
  not NOT_11544(II36981,g28074);
  not NOT_11545(g28244,II36981);
  not NOT_11546(II36984,g28013);
  not NOT_11547(g28245,II36984);
  not NOT_11548(II36987,g28033);
  not NOT_11549(g28246,II36987);
  not NOT_11550(II36990,g28054);
  not NOT_11551(g28247,II36990);
  not NOT_11552(II36993,g28034);
  not NOT_11553(g28248,II36993);
  not NOT_11554(II36996,g28055);
  not NOT_11555(g28249,II36996);
  not NOT_11556(II36999,g28076);
  not NOT_11557(g28250,II36999);
  not NOT_11558(II37002,g28056);
  not NOT_11559(g28251,II37002);
  not NOT_11560(II37005,g28077);
  not NOT_11561(g28252,II37005);
  not NOT_11562(II37008,g28096);
  not NOT_11563(g28253,II37008);
  not NOT_11564(II37011,g28078);
  not NOT_11565(g28254,II37011);
  not NOT_11566(II37014,g28097);
  not NOT_11567(g28255,II37014);
  not NOT_11568(II37017,g28113);
  not NOT_11569(g28256,II37017);
  not NOT_11570(II37020,g27910);
  not NOT_11571(g28257,II37020);
  not NOT_11572(II37023,g27799);
  not NOT_11573(g28258,II37023);
  not NOT_11574(II37026,g27998);
  not NOT_11575(g28259,II37026);
  not NOT_11576(II37029,g28016);
  not NOT_11577(g28260,II37029);
  not NOT_11578(II37032,g28037);
  not NOT_11579(g28261,II37032);
  not NOT_11580(II37035,g28017);
  not NOT_11581(g28262,II37035);
  not NOT_11582(II37038,g28038);
  not NOT_11583(g28263,II37038);
  not NOT_11584(II37041,g28060);
  not NOT_11585(g28264,II37041);
  not NOT_11586(II37044,g28039);
  not NOT_11587(g28265,II37044);
  not NOT_11588(II37047,g28061);
  not NOT_11589(g28266,II37047);
  not NOT_11590(II37050,g28081);
  not NOT_11591(g28267,II37050);
  not NOT_11592(II37053,g28062);
  not NOT_11593(g28268,II37053);
  not NOT_11594(II37056,g28082);
  not NOT_11595(g28269,II37056);
  not NOT_11596(II37059,g28099);
  not NOT_11597(g28270,II37059);
  not NOT_11598(II37062,g28040);
  not NOT_11599(g28271,II37062);
  not NOT_11600(II37065,g28063);
  not NOT_11601(g28272,II37065);
  not NOT_11602(II37068,g28083);
  not NOT_11603(g28273,II37068);
  not NOT_11604(II37071,g28064);
  not NOT_11605(g28274,II37071);
  not NOT_11606(II37074,g28084);
  not NOT_11607(g28275,II37074);
  not NOT_11608(II37077,g28101);
  not NOT_11609(g28276,II37077);
  not NOT_11610(II37080,g28085);
  not NOT_11611(g28277,II37080);
  not NOT_11612(II37083,g28102);
  not NOT_11613(g28278,II37083);
  not NOT_11614(II37086,g28114);
  not NOT_11615(g28279,II37086);
  not NOT_11616(II37089,g28103);
  not NOT_11617(g28280,II37089);
  not NOT_11618(II37092,g28115);
  not NOT_11619(g28281,II37092);
  not NOT_11620(II37095,g28124);
  not NOT_11621(g28282,II37095);
  not NOT_11622(II37098,g27918);
  not NOT_11623(g28283,II37098);
  not NOT_11624(II37101,g27805);
  not NOT_11625(g28284,II37101);
  not NOT_11626(II37104,g28021);
  not NOT_11627(g28285,II37104);
  not NOT_11628(II37107,g28043);
  not NOT_11629(g28286,II37107);
  not NOT_11630(II37110,g28067);
  not NOT_11631(g28287,II37110);
  not NOT_11632(II37113,g28044);
  not NOT_11633(g28288,II37113);
  not NOT_11634(II37116,g28068);
  not NOT_11635(g28289,II37116);
  not NOT_11636(II37119,g28089);
  not NOT_11637(g28290,II37119);
  not NOT_11638(II37122,g28069);
  not NOT_11639(g28291,II37122);
  not NOT_11640(II37125,g28090);
  not NOT_11641(g28292,II37125);
  not NOT_11642(II37128,g28106);
  not NOT_11643(g28293,II37128);
  not NOT_11644(II37131,g28091);
  not NOT_11645(g28294,II37131);
  not NOT_11646(II37134,g28107);
  not NOT_11647(g28295,II37134);
  not NOT_11648(II37137,g28117);
  not NOT_11649(g28296,II37137);
  not NOT_11650(II37140,g28070);
  not NOT_11651(g28297,II37140);
  not NOT_11652(II37143,g28092);
  not NOT_11653(g28298,II37143);
  not NOT_11654(II37146,g28108);
  not NOT_11655(g28299,II37146);
  not NOT_11656(II37149,g28093);
  not NOT_11657(g28300,II37149);
  not NOT_11658(II37152,g28109);
  not NOT_11659(g28301,II37152);
  not NOT_11660(II37155,g28119);
  not NOT_11661(g28302,II37155);
  not NOT_11662(II37158,g28110);
  not NOT_11663(g28303,II37158);
  not NOT_11664(II37161,g28120);
  not NOT_11665(g28304,II37161);
  not NOT_11666(II37164,g28125);
  not NOT_11667(g28305,II37164);
  not NOT_11668(II37167,g28121);
  not NOT_11669(g28306,II37167);
  not NOT_11670(II37170,g28126);
  not NOT_11671(g28307,II37170);
  not NOT_11672(II37173,g28132);
  not NOT_11673(g28308,II37173);
  not NOT_11674(II37176,g27927);
  not NOT_11675(g28309,II37176);
  not NOT_11676(II37179,g27784);
  not NOT_11677(g28310,II37179);
  not NOT_11678(II37182,g27791);
  not NOT_11679(g28311,II37182);
  not NOT_11680(II37185,g27797);
  not NOT_11681(g28312,II37185);
  not NOT_11682(II37188,g27785);
  not NOT_11683(g28313,II37188);
  not NOT_11684(II37191,g27792);
  not NOT_11685(g28314,II37191);
  not NOT_11686(II37194,g27800);
  not NOT_11687(g28315,II37194);
  not NOT_11688(II37197,g27903);
  not NOT_11689(g28316,II37197);
  not NOT_11690(II37200,g27907);
  not NOT_11691(g28317,II37200);
  not NOT_11692(II37203,g27912);
  not NOT_11693(g28318,II37203);
  not NOT_11694(II37228,g28194);
  not NOT_11695(g28341,II37228);
  not NOT_11696(II37232,g28200);
  not NOT_11697(g28343,II37232);
  not NOT_11698(II37238,g28179);
  not NOT_11699(g28347,II37238);
  not NOT_11700(II37252,g28200);
  not NOT_11701(g28359,II37252);
  not NOT_11702(II37260,g28179);
  not NOT_11703(g28365,II37260);
  not NOT_11704(II37266,g28200);
  not NOT_11705(g28369,II37266);
  not NOT_11706(II37269,g28145);
  not NOT_11707(g28370,II37269);
  not NOT_11708(II37273,g28179);
  not NOT_11709(g28372,II37273);
  not NOT_11710(II37277,g28146);
  not NOT_11711(g28374,II37277);
  not NOT_11712(II37280,g28179);
  not NOT_11713(g28375,II37280);
  not NOT_11714(II37284,g28147);
  not NOT_11715(g28377,II37284);
  not NOT_11716(II37291,g28148);
  not NOT_11717(g28382,II37291);
  not NOT_11718(II37319,g28149);
  not NOT_11719(g28390,II37319);
  not NOT_11720(II37330,g28194);
  not NOT_11721(g28393,II37330);
  not NOT_11722(II37334,g28194);
  not NOT_11723(g28395,II37334);
  not NOT_11724(g28419,g28151);
  not NOT_11725(II37379,g28199);
  not NOT_11726(g28432,II37379);
  not NOT_11727(II37386,g28194);
  not NOT_11728(g28437,II37386);
  not NOT_11729(II37394,g27718);
  not NOT_11730(g28443,II37394);
  not NOT_11731(II37400,g28200);
  not NOT_11732(g28447,II37400);
  not NOT_11733(II37410,g27722);
  not NOT_11734(g28455,II37410);
  not NOT_11735(II37415,g28179);
  not NOT_11736(g28458,II37415);
  not NOT_11737(II37426,g27724);
  not NOT_11738(g28467,II37426);
  not NOT_11739(g28483,g27776);
  not NOT_11740(g28491,g27780);
  not NOT_11741(g28496,g27787);
  not NOT_11742(II37459,g27759);
  not NOT_11743(g28498,II37459);
  not NOT_11744(g28500,g27794);
  not NOT_11745(II37467,g27760);
  not NOT_11746(g28524,II37467);
  not NOT_11747(II37471,g27761);
  not NOT_11748(g28526,II37471);
  not NOT_11749(II37474,g27762);
  not NOT_11750(g28527,II37474);
  not NOT_11751(II37481,g27763);
  not NOT_11752(g28552,II37481);
  not NOT_11753(II37484,g27764);
  not NOT_11754(g28553,II37484);
  not NOT_11755(g28554,g27806);
  not NOT_11756(II37488,g27765);
  not NOT_11757(g28555,II37488);
  not NOT_11758(II37494,g27766);
  not NOT_11759(g28579,II37494);
  not NOT_11760(II37497,g27767);
  not NOT_11761(g28580,II37497);
  not NOT_11762(g28581,g27817);
  not NOT_11763(g28582,g27820);
  not NOT_11764(II37502,g27768);
  not NOT_11765(g28583,II37502);
  not NOT_11766(II37508,g27769);
  not NOT_11767(g28607,II37508);
  not NOT_11768(g28608,g27831);
  not NOT_11769(g28609,g27839);
  not NOT_11770(g28610,g27843);
  not NOT_11771(II37514,g27771);
  not NOT_11772(g28611,II37514);
  not NOT_11773(g28612,g28046);
  not NOT_11774(g28616,g27847);
  not NOT_11775(g28617,g27858);
  not NOT_11776(g28618,g27861);
  not NOT_11777(g28619,g28075);
  not NOT_11778(g28623,g27872);
  not NOT_11779(g28624,g27879);
  not NOT_11780(g28625,g28100);
  not NOT_11781(g28629,g27889);
  not NOT_11782(g28630,g28118);
  not NOT_11783(g28638,g28200);
  not NOT_11784(g28639,g27919);
  not NOT_11785(g28640,g27928);
  not NOT_11786(g28641,g27932);
  not NOT_11787(g28642,g27939);
  not NOT_11788(g28643,g27942);
  not NOT_11789(g28644,g27946);
  not NOT_11790(g28645,g27952);
  not NOT_11791(g28646,g27956);
  not NOT_11792(g28647,g27959);
  not NOT_11793(g28648,g27965);
  not NOT_11794(g28649,g27973);
  not NOT_11795(g28650,g27977);
  not NOT_11796(g28651,g27981);
  not NOT_11797(g28652,g27994);
  not NOT_11798(g28653,g27999);
  not NOT_11799(g28655,g28018);
  not NOT_11800(II37566,g28370);
  not NOT_11801(g28673,II37566);
  not NOT_11802(II37569,g28498);
  not NOT_11803(g28674,II37569);
  not NOT_11804(II37572,g28524);
  not NOT_11805(g28675,II37572);
  not NOT_11806(II37575,g28527);
  not NOT_11807(g28676,II37575);
  not NOT_11808(II37578,g28432);
  not NOT_11809(g28677,II37578);
  not NOT_11810(II37581,g28374);
  not NOT_11811(g28678,II37581);
  not NOT_11812(II37584,g28526);
  not NOT_11813(g28679,II37584);
  not NOT_11814(II37587,g28552);
  not NOT_11815(g28680,II37587);
  not NOT_11816(II37590,g28555);
  not NOT_11817(g28681,II37590);
  not NOT_11818(II37593,g28443);
  not NOT_11819(g28682,II37593);
  not NOT_11820(II37596,g28377);
  not NOT_11821(g28683,II37596);
  not NOT_11822(II37599,g28553);
  not NOT_11823(g28684,II37599);
  not NOT_11824(II37602,g28579);
  not NOT_11825(g28685,II37602);
  not NOT_11826(II37605,g28583);
  not NOT_11827(g28686,II37605);
  not NOT_11828(II37608,g28455);
  not NOT_11829(g28687,II37608);
  not NOT_11830(II37611,g28382);
  not NOT_11831(g28688,II37611);
  not NOT_11832(II37614,g28580);
  not NOT_11833(g28689,II37614);
  not NOT_11834(II37617,g28607);
  not NOT_11835(g28690,II37617);
  not NOT_11836(II37620,g28611);
  not NOT_11837(g28691,II37620);
  not NOT_11838(II37623,g28467);
  not NOT_11839(g28692,II37623);
  not NOT_11840(II37626,g28393);
  not NOT_11841(g28693,II37626);
  not NOT_11842(II37629,g28369);
  not NOT_11843(g28694,II37629);
  not NOT_11844(II37632,g28372);
  not NOT_11845(g28695,II37632);
  not NOT_11846(II37635,g28390);
  not NOT_11847(g28696,II37635);
  not NOT_11848(II37638,g28395);
  not NOT_11849(g28697,II37638);
  not NOT_11850(II37641,g28375);
  not NOT_11851(g28698,II37641);
  not NOT_11852(II37644,g28341);
  not NOT_11853(g28699,II37644);
  not NOT_11854(II37647,g28343);
  not NOT_11855(g28700,II37647);
  not NOT_11856(II37650,g28347);
  not NOT_11857(g28701,II37650);
  not NOT_11858(II37653,g28359);
  not NOT_11859(g28702,II37653);
  not NOT_11860(II37656,g28365);
  not NOT_11861(g28703,II37656);
  not NOT_11862(II37659,g28437);
  not NOT_11863(g28704,II37659);
  not NOT_11864(II37662,g28447);
  not NOT_11865(g28705,II37662);
  not NOT_11866(II37665,g28458);
  not NOT_11867(g28706,II37665);
  not NOT_11868(g28720,g28495);
  not NOT_11869(g28721,g28490);
  not NOT_11870(g28723,g28528);
  not NOT_11871(g28725,g28499);
  not NOT_11872(g28727,g28489);
  not NOT_11873(g28730,g28470);
  not NOT_11874(g28734,g28525);
  not NOT_11875(g28740,g28488);
  not NOT_11876(II37702,g28512);
  not NOT_11877(g28741,II37702);
  not NOT_11878(II37712,g28512);
  not NOT_11879(g28751,II37712);
  not NOT_11880(II37716,g28540);
  not NOT_11881(g28755,II37716);
  not NOT_11882(II37725,g28540);
  not NOT_11883(g28764,II37725);
  not NOT_11884(II37729,g28567);
  not NOT_11885(g28768,II37729);
  not NOT_11886(II37736,g28567);
  not NOT_11887(g28775,II37736);
  not NOT_11888(II37740,g28595);
  not NOT_11889(g28779,II37740);
  not NOT_11890(II37746,g28595);
  not NOT_11891(g28785,II37746);
  not NOT_11892(II37752,g28512);
  not NOT_11893(g28791,II37752);
  not NOT_11894(II37757,g28512);
  not NOT_11895(g28796,II37757);
  not NOT_11896(II37760,g28540);
  not NOT_11897(g28799,II37760);
  not NOT_11898(II37765,g28512);
  not NOT_11899(g28804,II37765);
  not NOT_11900(II37768,g28540);
  not NOT_11901(g28807,II37768);
  not NOT_11902(II37771,g28567);
  not NOT_11903(g28810,II37771);
  not NOT_11904(II37775,g28540);
  not NOT_11905(g28814,II37775);
  not NOT_11906(II37778,g28567);
  not NOT_11907(g28817,II37778);
  not NOT_11908(II37781,g28595);
  not NOT_11909(g28820,II37781);
  not NOT_11910(II37784,g28567);
  not NOT_11911(g28823,II37784);
  not NOT_11912(II37787,g28595);
  not NOT_11913(g28826,II37787);
  not NOT_11914(II37790,g28595);
  not NOT_11915(g28829,II37790);
  not NOT_11916(II37793,g28638);
  not NOT_11917(g28832,II37793);
  not NOT_11918(II37796,g28634);
  not NOT_11919(g28833,II37796);
  not NOT_11920(II37800,g28635);
  not NOT_11921(g28835,II37800);
  not NOT_11922(II37804,g28636);
  not NOT_11923(g28837,II37804);
  not NOT_11924(II37808,g28637);
  not NOT_11925(g28839,II37808);
  not NOT_11926(g28855,g28409);
  not NOT_11927(g28859,g28413);
  not NOT_11928(g28863,g28417);
  not NOT_11929(g28867,g28418);
  not NOT_11930(II37842,g28501);
  not NOT_11931(g28871,II37842);
  not NOT_11932(II37846,g28501);
  not NOT_11933(g28877,II37846);
  not NOT_11934(II37851,g28668);
  not NOT_11935(g28882,II37851);
  not NOT_11936(II37854,g28529);
  not NOT_11937(g28883,II37854);
  not NOT_11938(II37858,g28501);
  not NOT_11939(g28889,II37858);
  not NOT_11940(II37863,g28529);
  not NOT_11941(g28894,II37863);
  not NOT_11942(II37868,g28321);
  not NOT_11943(g28899,II37868);
  not NOT_11944(II37871,g28556);
  not NOT_11945(g28900,II37871);
  not NOT_11946(II37875,g28501);
  not NOT_11947(g28906,II37875);
  not NOT_11948(II37880,g28529);
  not NOT_11949(g28911,II37880);
  not NOT_11950(II37885,g28556);
  not NOT_11951(g28916,II37885);
  not NOT_11952(II37891,g28325);
  not NOT_11953(g28924,II37891);
  not NOT_11954(II37894,g28584);
  not NOT_11955(g28925,II37894);
  not NOT_11956(II37897,g28501);
  not NOT_11957(g28928,II37897);
  not NOT_11958(II37901,g28529);
  not NOT_11959(g28932,II37901);
  not NOT_11960(II37906,g28556);
  not NOT_11961(g28937,II37906);
  not NOT_11962(II37912,g28584);
  not NOT_11963(g28945,II37912);
  not NOT_11964(II37917,g28328);
  not NOT_11965(g28950,II37917);
  not NOT_11966(II37920,g28501);
  not NOT_11967(g28951,II37920);
  not NOT_11968(II37924,g28529);
  not NOT_11969(g28955,II37924);
  not NOT_11970(II37928,g28556);
  not NOT_11971(g28959,II37928);
  not NOT_11972(II37934,g28584);
  not NOT_11973(g28967,II37934);
  not NOT_11974(II37939,g28501);
  not NOT_11975(g28972,II37939);
  not NOT_11976(II37942,g28501);
  not NOT_11977(g28975,II37942);
  not NOT_11978(II37946,g28529);
  not NOT_11979(g28979,II37946);
  not NOT_11980(II37950,g28556);
  not NOT_11981(g28983,II37950);
  not NOT_11982(II37956,g28584);
  not NOT_11983(g28993,II37956);
  not NOT_11984(II37961,g28501);
  not NOT_11985(g28998,II37961);
  not NOT_11986(II37965,g28529);
  not NOT_11987(g29002,II37965);
  not NOT_11988(II37968,g28529);
  not NOT_11989(g29005,II37968);
  not NOT_11990(II37973,g28556);
  not NOT_11991(g29010,II37973);
  not NOT_11992(II37978,g28584);
  not NOT_11993(g29019,II37978);
  not NOT_11994(II37982,g28501);
  not NOT_11995(g29023,II37982);
  not NOT_11996(II37986,g28529);
  not NOT_11997(g29027,II37986);
  not NOT_11998(II37991,g28556);
  not NOT_11999(g29032,II37991);
  not NOT_12000(II37994,g28556);
  not NOT_12001(g29035,II37994);
  not NOT_12002(II37999,g28584);
  not NOT_12003(g29042,II37999);
  not NOT_12004(II38003,g28529);
  not NOT_12005(g29046,II38003);
  not NOT_12006(II38007,g28556);
  not NOT_12007(g29050,II38007);
  not NOT_12008(II38011,g28584);
  not NOT_12009(g29054,II38011);
  not NOT_12010(II38014,g28584);
  not NOT_12011(g29057,II38014);
  not NOT_12012(II38018,g28342);
  not NOT_12013(g29061,II38018);
  not NOT_12014(II38024,g28556);
  not NOT_12015(g29065,II38024);
  not NOT_12016(II38028,g28584);
  not NOT_12017(g29069,II38028);
  not NOT_12018(II38032,g28344);
  not NOT_12019(g29073,II38032);
  not NOT_12020(II38035,g28345);
  not NOT_12021(g29074,II38035);
  not NOT_12022(II38038,g28346);
  not NOT_12023(g29075,II38038);
  not NOT_12024(II38042,g28584);
  not NOT_12025(g29077,II38042);
  not NOT_12026(II38046,g28348);
  not NOT_12027(g29081,II38046);
  not NOT_12028(II38049,g28349);
  not NOT_12029(g29082,II38049);
  not NOT_12030(II38053,g28350);
  not NOT_12031(g29084,II38053);
  not NOT_12032(II38056,g28351);
  not NOT_12033(g29085,II38056);
  not NOT_12034(II38059,g28352);
  not NOT_12035(g29086,II38059);
  not NOT_12036(II38064,g28353);
  not NOT_12037(g29089,II38064);
  not NOT_12038(II38068,g28354);
  not NOT_12039(g29091,II38068);
  not NOT_12040(II38071,g28355);
  not NOT_12041(g29092,II38071);
  not NOT_12042(II38074,g28356);
  not NOT_12043(g29093,II38074);
  not NOT_12044(II38077,g28357);
  not NOT_12045(g29094,II38077);
  not NOT_12046(II38080,g28358);
  not NOT_12047(g29095,II38080);
  not NOT_12048(II38085,g28360);
  not NOT_12049(g29098,II38085);
  not NOT_12050(II38088,g28361);
  not NOT_12051(g29099,II38088);
  not NOT_12052(II38091,g28362);
  not NOT_12053(g29100,II38091);
  not NOT_12054(II38094,g28363);
  not NOT_12055(g29101,II38094);
  not NOT_12056(II38097,g28364);
  not NOT_12057(g29102,II38097);
  not NOT_12058(II38101,g28366);
  not NOT_12059(g29104,II38101);
  not NOT_12060(II38104,g28367);
  not NOT_12061(g29105,II38104);
  not NOT_12062(II38107,g28368);
  not NOT_12063(g29106,II38107);
  not NOT_12064(II38111,g28371);
  not NOT_12065(g29108,II38111);
  not NOT_12066(II38119,g28420);
  not NOT_12067(g29117,II38119);
  not NOT_12068(II38122,g28421);
  not NOT_12069(g29118,II38122);
  not NOT_12070(II38125,g28425);
  not NOT_12071(g29119,II38125);
  not NOT_12072(II38128,g28419);
  not NOT_12073(g29120,II38128);
  not NOT_12074(II38136,g28833);
  not NOT_12075(g29131,II38136);
  not NOT_12076(II38139,g29061);
  not NOT_12077(g29132,II38139);
  not NOT_12078(II38142,g29073);
  not NOT_12079(g29133,II38142);
  not NOT_12080(II38145,g29081);
  not NOT_12081(g29134,II38145);
  not NOT_12082(II38148,g29074);
  not NOT_12083(g29135,II38148);
  not NOT_12084(II38151,g29082);
  not NOT_12085(g29136,II38151);
  not NOT_12086(II38154,g29089);
  not NOT_12087(g29137,II38154);
  not NOT_12088(II38157,g28882);
  not NOT_12089(g29138,II38157);
  not NOT_12090(II38160,g28835);
  not NOT_12091(g29139,II38160);
  not NOT_12092(II38163,g29075);
  not NOT_12093(g29140,II38163);
  not NOT_12094(II38166,g29084);
  not NOT_12095(g29141,II38166);
  not NOT_12096(II38169,g29091);
  not NOT_12097(g29142,II38169);
  not NOT_12098(II38172,g29085);
  not NOT_12099(g29143,II38172);
  not NOT_12100(II38175,g29092);
  not NOT_12101(g29144,II38175);
  not NOT_12102(II38178,g29098);
  not NOT_12103(g29145,II38178);
  not NOT_12104(II38181,g28899);
  not NOT_12105(g29146,II38181);
  not NOT_12106(II38184,g28837);
  not NOT_12107(g29147,II38184);
  not NOT_12108(II38187,g29086);
  not NOT_12109(g29148,II38187);
  not NOT_12110(II38190,g29093);
  not NOT_12111(g29149,II38190);
  not NOT_12112(II38193,g29099);
  not NOT_12113(g29150,II38193);
  not NOT_12114(II38196,g29094);
  not NOT_12115(g29151,II38196);
  not NOT_12116(II38199,g29100);
  not NOT_12117(g29152,II38199);
  not NOT_12118(II38202,g29104);
  not NOT_12119(g29153,II38202);
  not NOT_12120(II38205,g28924);
  not NOT_12121(g29154,II38205);
  not NOT_12122(II38208,g28839);
  not NOT_12123(g29155,II38208);
  not NOT_12124(II38211,g29095);
  not NOT_12125(g29156,II38211);
  not NOT_12126(II38214,g29101);
  not NOT_12127(g29157,II38214);
  not NOT_12128(II38217,g29105);
  not NOT_12129(g29158,II38217);
  not NOT_12130(II38220,g29102);
  not NOT_12131(g29159,II38220);
  not NOT_12132(II38223,g29106);
  not NOT_12133(g29160,II38223);
  not NOT_12134(II38226,g29108);
  not NOT_12135(g29161,II38226);
  not NOT_12136(II38229,g28950);
  not NOT_12137(g29162,II38229);
  not NOT_12138(II38232,g29117);
  not NOT_12139(g29163,II38232);
  not NOT_12140(II38235,g29118);
  not NOT_12141(g29164,II38235);
  not NOT_12142(II38238,g29119);
  not NOT_12143(g29165,II38238);
  not NOT_12144(II38241,g28832);
  not NOT_12145(g29166,II38241);
  not NOT_12146(II38245,g28920);
  not NOT_12147(g29168,II38245);
  not NOT_12148(II38250,g28941);
  not NOT_12149(g29171,II38250);
  not NOT_12150(II38258,g28963);
  not NOT_12151(g29177,II38258);
  not NOT_12152(II38272,g29013);
  not NOT_12153(g29189,II38272);
  not NOT_12154(II38275,g28987);
  not NOT_12155(g29190,II38275);
  not NOT_12156(II38278,g28963);
  not NOT_12157(g29191,II38278);
  not NOT_12158(g29192,g28954);
  not NOT_12159(II38282,g28941);
  not NOT_12160(g29193,II38282);
  not NOT_12161(II38321,g29113);
  not NOT_12162(g29230,II38321);
  not NOT_12163(II38330,g29120);
  not NOT_12164(g29237,II38330);
  not NOT_12165(II38339,g29120);
  not NOT_12166(g29244,II38339);
  not NOT_12167(II38342,g28886);
  not NOT_12168(g29245,II38342);
  not NOT_12169(II38345,g29109);
  not NOT_12170(g29246,II38345);
  not NOT_12171(II38348,g28874);
  not NOT_12172(g29247,II38348);
  not NOT_12173(II38352,g29110);
  not NOT_12174(g29249,II38352);
  not NOT_12175(II38355,g29039);
  not NOT_12176(g29250,II38355);
  not NOT_12177(II38360,g29111);
  not NOT_12178(g29253,II38360);
  not NOT_12179(II38363,g29016);
  not NOT_12180(g29254,II38363);
  not NOT_12181(II38369,g29112);
  not NOT_12182(g29258,II38369);
  not NOT_12183(g29266,g28741);
  not NOT_12184(II38386,g28734);
  not NOT_12185(g29267,II38386);
  not NOT_12186(g29268,g28751);
  not NOT_12187(g29269,g28755);
  not NOT_12188(II38391,g28730);
  not NOT_12189(g29270,II38391);
  not NOT_12190(g29271,g28764);
  not NOT_12191(g29272,g28768);
  not NOT_12192(II38396,g28727);
  not NOT_12193(g29273,II38396);
  not NOT_12194(g29274,g28775);
  not NOT_12195(g29275,g28779);
  not NOT_12196(II38401,g28725);
  not NOT_12197(g29276,II38401);
  not NOT_12198(g29277,g28785);
  not NOT_12199(II38405,g28723);
  not NOT_12200(g29278,II38405);
  not NOT_12201(II38408,g28721);
  not NOT_12202(g29279,II38408);
  not NOT_12203(g29280,g28791);
  not NOT_12204(II38412,g28720);
  not NOT_12205(g29281,II38412);
  not NOT_12206(g29282,g28796);
  not NOT_12207(g29283,g28799);
  not NOT_12208(g29285,g28804);
  not NOT_12209(g29286,g28807);
  not NOT_12210(g29287,g28810);
  not NOT_12211(II38421,g28740);
  not NOT_12212(g29288,II38421);
  not NOT_12213(g29290,g28814);
  not NOT_12214(g29291,g28817);
  not NOT_12215(g29292,g28820);
  not NOT_12216(II38428,g28732);
  not NOT_12217(g29293,II38428);
  not NOT_12218(g29295,g28823);
  not NOT_12219(g29296,g28826);
  not NOT_12220(II38434,g28735);
  not NOT_12221(g29297,II38434);
  not NOT_12222(II38437,g28736);
  not NOT_12223(g29298,II38437);
  not NOT_12224(II38440,g28738);
  not NOT_12225(g29299,II38440);
  not NOT_12226(g29301,g28829);
  not NOT_12227(II38447,g28744);
  not NOT_12228(g29304,II38447);
  not NOT_12229(II38450,g28745);
  not NOT_12230(g29305,II38450);
  not NOT_12231(II38453,g28746);
  not NOT_12232(g29306,II38453);
  not NOT_12233(II38456,g28747);
  not NOT_12234(g29307,II38456);
  not NOT_12235(II38459,g28749);
  not NOT_12236(g29308,II38459);
  not NOT_12237(II38462,g29120);
  not NOT_12238(g29309,II38462);
  not NOT_12239(II38466,g28754);
  not NOT_12240(g29311,II38466);
  not NOT_12241(II38471,g28758);
  not NOT_12242(g29314,II38471);
  not NOT_12243(II38474,g28759);
  not NOT_12244(g29315,II38474);
  not NOT_12245(II38477,g28760);
  not NOT_12246(g29316,II38477);
  not NOT_12247(II38480,g28761);
  not NOT_12248(g29317,II38480);
  not NOT_12249(II38483,g28990);
  not NOT_12250(g29318,II38483);
  not NOT_12251(II38486,g28763);
  not NOT_12252(g29319,II38486);
  not NOT_12253(II38491,g28767);
  not NOT_12254(g29322,II38491);
  not NOT_12255(II38496,g28771);
  not NOT_12256(g29325,II38496);
  not NOT_12257(II38499,g28772);
  not NOT_12258(g29326,II38499);
  not NOT_12259(II38502,g28773);
  not NOT_12260(g29327,II38502);
  not NOT_12261(II38505,g28774);
  not NOT_12262(g29328,II38505);
  not NOT_12263(II38510,g28778);
  not NOT_12264(g29331,II38510);
  not NOT_12265(II38515,g28782);
  not NOT_12266(g29334,II38515);
  not NOT_12267(II38518,g28783);
  not NOT_12268(g29335,II38518);
  not NOT_12269(II38524,g28788);
  not NOT_12270(g29339,II38524);
  not NOT_12271(II38536,g28920);
  not NOT_12272(g29349,II38536);
  not NOT_12273(II38539,g29113);
  not NOT_12274(g29350,II38539);
  not NOT_12275(g29356,g29120);
  not NOT_12276(g29358,g29120);
  not NOT_12277(II38548,g28903);
  not NOT_12278(g29359,II38548);
  not NOT_12279(g29360,g28871);
  not NOT_12280(g29361,g28877);
  not NOT_12281(g29362,g28883);
  not NOT_12282(g29363,g28889);
  not NOT_12283(g29364,g28894);
  not NOT_12284(g29365,g28900);
  not NOT_12285(g29366,g28906);
  not NOT_12286(g29367,g28911);
  not NOT_12287(g29368,g28916);
  not NOT_12288(g29369,g28925);
  not NOT_12289(g29370,g28928);
  not NOT_12290(g29371,g28932);
  not NOT_12291(g29372,g28937);
  not NOT_12292(g29373,g28945);
  not NOT_12293(g29374,g28951);
  not NOT_12294(g29375,g28955);
  not NOT_12295(g29376,g28959);
  not NOT_12296(g29377,g28967);
  not NOT_12297(g29378,g28972);
  not NOT_12298(g29379,g28975);
  not NOT_12299(g29380,g28979);
  not NOT_12300(g29381,g28983);
  not NOT_12301(g29382,g28993);
  not NOT_12302(g29383,g28998);
  not NOT_12303(g29384,g29002);
  not NOT_12304(g29385,g29005);
  not NOT_12305(g29386,g29010);
  not NOT_12306(g29387,g29019);
  not NOT_12307(g29388,g29023);
  not NOT_12308(g29389,g29027);
  not NOT_12309(g29390,g29032);
  not NOT_12310(g29391,g29035);
  not NOT_12311(g29392,g29042);
  not NOT_12312(g29393,g29046);
  not NOT_12313(g29394,g29050);
  not NOT_12314(g29395,g29054);
  not NOT_12315(g29396,g29057);
  not NOT_12316(g29397,g29065);
  not NOT_12317(g29398,g29069);
  not NOT_12318(II38591,g28987);
  not NOT_12319(g29400,II38591);
  not NOT_12320(II38594,g28990);
  not NOT_12321(g29401,II38594);
  not NOT_12322(g29402,g29077);
  not NOT_12323(II38599,g29013);
  not NOT_12324(g29404,II38599);
  not NOT_12325(II38602,g29016);
  not NOT_12326(g29405,II38602);
  not NOT_12327(II38606,g29039);
  not NOT_12328(g29407,II38606);
  not NOT_12329(II38609,g28874);
  not NOT_12330(g29408,II38609);
  not NOT_12331(II38613,g28886);
  not NOT_12332(g29410,II38613);
  not NOT_12333(II38617,g28903);
  not NOT_12334(g29412,II38617);
  not NOT_12335(II38620,g29246);
  not NOT_12336(g29413,II38620);
  not NOT_12337(II38623,g29293);
  not NOT_12338(g29414,II38623);
  not NOT_12339(II38626,g29297);
  not NOT_12340(g29415,II38626);
  not NOT_12341(II38629,g29304);
  not NOT_12342(g29416,II38629);
  not NOT_12343(II38632,g29298);
  not NOT_12344(g29417,II38632);
  not NOT_12345(II38635,g29305);
  not NOT_12346(g29418,II38635);
  not NOT_12347(II38638,g29311);
  not NOT_12348(g29419,II38638);
  not NOT_12349(II38641,g29249);
  not NOT_12350(g29420,II38641);
  not NOT_12351(II38644,g29299);
  not NOT_12352(g29421,II38644);
  not NOT_12353(II38647,g29306);
  not NOT_12354(g29422,II38647);
  not NOT_12355(II38650,g29314);
  not NOT_12356(g29423,II38650);
  not NOT_12357(II38653,g29307);
  not NOT_12358(g29424,II38653);
  not NOT_12359(II38656,g29315);
  not NOT_12360(g29425,II38656);
  not NOT_12361(II38659,g29322);
  not NOT_12362(g29426,II38659);
  not NOT_12363(II38662,g29253);
  not NOT_12364(g29427,II38662);
  not NOT_12365(II38665,g29412);
  not NOT_12366(g29428,II38665);
  not NOT_12367(II38668,g29168);
  not NOT_12368(g29429,II38668);
  not NOT_12369(II38671,g29171);
  not NOT_12370(g29430,II38671);
  not NOT_12371(II38674,g29177);
  not NOT_12372(g29431,II38674);
  not NOT_12373(II38677,g29400);
  not NOT_12374(g29432,II38677);
  not NOT_12375(II38680,g29404);
  not NOT_12376(g29433,II38680);
  not NOT_12377(II38683,g29308);
  not NOT_12378(g29434,II38683);
  not NOT_12379(II38686,g29316);
  not NOT_12380(g29435,II38686);
  not NOT_12381(II38689,g29325);
  not NOT_12382(g29436,II38689);
  not NOT_12383(II38692,g29317);
  not NOT_12384(g29437,II38692);
  not NOT_12385(II38695,g29326);
  not NOT_12386(g29438,II38695);
  not NOT_12387(II38698,g29331);
  not NOT_12388(g29439,II38698);
  not NOT_12389(II38701,g29401);
  not NOT_12390(g29440,II38701);
  not NOT_12391(II38704,g29405);
  not NOT_12392(g29441,II38704);
  not NOT_12393(II38707,g29407);
  not NOT_12394(g29442,II38707);
  not NOT_12395(II38710,g29408);
  not NOT_12396(g29443,II38710);
  not NOT_12397(II38713,g29410);
  not NOT_12398(g29444,II38713);
  not NOT_12399(II38716,g29230);
  not NOT_12400(g29445,II38716);
  not NOT_12401(II38719,g29258);
  not NOT_12402(g29446,II38719);
  not NOT_12403(II38722,g29319);
  not NOT_12404(g29447,II38722);
  not NOT_12405(II38725,g29327);
  not NOT_12406(g29448,II38725);
  not NOT_12407(II38728,g29334);
  not NOT_12408(g29449,II38728);
  not NOT_12409(II38731,g29328);
  not NOT_12410(g29450,II38731);
  not NOT_12411(II38734,g29335);
  not NOT_12412(g29451,II38734);
  not NOT_12413(II38737,g29339);
  not NOT_12414(g29452,II38737);
  not NOT_12415(II38740,g29288);
  not NOT_12416(g29453,II38740);
  not NOT_12417(II38743,g29267);
  not NOT_12418(g29454,II38743);
  not NOT_12419(II38746,g29270);
  not NOT_12420(g29455,II38746);
  not NOT_12421(II38749,g29273);
  not NOT_12422(g29456,II38749);
  not NOT_12423(II38752,g29276);
  not NOT_12424(g29457,II38752);
  not NOT_12425(II38755,g29278);
  not NOT_12426(g29458,II38755);
  not NOT_12427(II38758,g29279);
  not NOT_12428(g29459,II38758);
  not NOT_12429(II38761,g29281);
  not NOT_12430(g29460,II38761);
  not NOT_12431(II38764,g29237);
  not NOT_12432(g29461,II38764);
  not NOT_12433(II38767,g29244);
  not NOT_12434(g29462,II38767);
  not NOT_12435(II38770,g29309);
  not NOT_12436(g29463,II38770);
  not NOT_12437(g29491,g29350);
  not NOT_12438(II38801,g29358);
  not NOT_12439(g29495,II38801);
  not NOT_12440(II38804,g29353);
  not NOT_12441(g29496,II38804);
  not NOT_12442(II38807,g29356);
  not NOT_12443(g29497,II38807);
  not NOT_12444(II38817,g29354);
  not NOT_12445(g29499,II38817);
  not NOT_12446(II38827,g29355);
  not NOT_12447(g29501,II38827);
  not NOT_12448(II38838,g29357);
  not NOT_12449(g29504,II38838);
  not NOT_12450(II38848,g29167);
  not NOT_12451(g29506,II38848);
  not NOT_12452(II38851,g29169);
  not NOT_12453(g29507,II38851);
  not NOT_12454(II38854,g29170);
  not NOT_12455(g29508,II38854);
  not NOT_12456(II38857,g29172);
  not NOT_12457(g29509,II38857);
  not NOT_12458(II38860,g29173);
  not NOT_12459(g29510,II38860);
  not NOT_12460(II38863,g29178);
  not NOT_12461(g29511,II38863);
  not NOT_12462(II38866,g29179);
  not NOT_12463(g29512,II38866);
  not NOT_12464(II38869,g29181);
  not NOT_12465(g29513,II38869);
  not NOT_12466(II38872,g29182);
  not NOT_12467(g29514,II38872);
  not NOT_12468(II38875,g29184);
  not NOT_12469(g29515,II38875);
  not NOT_12470(II38878,g29185);
  not NOT_12471(g29516,II38878);
  not NOT_12472(II38881,g29187);
  not NOT_12473(g29517,II38881);
  not NOT_12474(II38885,g29192);
  not NOT_12475(g29519,II38885);
  not NOT_12476(II38898,g29194);
  not NOT_12477(g29530,II38898);
  not NOT_12478(II38905,g29197);
  not NOT_12479(g29535,II38905);
  not NOT_12480(II38909,g29198);
  not NOT_12481(g29537,II38909);
  not NOT_12482(II38916,g29201);
  not NOT_12483(g29542,II38916);
  not NOT_12484(II38920,g29204);
  not NOT_12485(g29544,II38920);
  not NOT_12486(II38924,g29205);
  not NOT_12487(g29546,II38924);
  not NOT_12488(II38931,g29209);
  not NOT_12489(g29551,II38931);
  not NOT_12490(II38936,g29212);
  not NOT_12491(g29554,II38936);
  not NOT_12492(II38940,g29213);
  not NOT_12493(g29556,II38940);
  not NOT_12494(II38947,g29218);
  not NOT_12495(g29561,II38947);
  not NOT_12496(II38951,g29221);
  not NOT_12497(g29563,II38951);
  not NOT_12498(II38958,g29226);
  not NOT_12499(g29568,II38958);
  not NOT_12500(II38975,g29348);
  not NOT_12501(g29583,II38975);
  not NOT_12502(II38999,g29496);
  not NOT_12503(g29627,II38999);
  not NOT_12504(II39002,g29506);
  not NOT_12505(g29628,II39002);
  not NOT_12506(II39005,g29507);
  not NOT_12507(g29629,II39005);
  not NOT_12508(II39008,g29509);
  not NOT_12509(g29630,II39008);
  not NOT_12510(II39011,g29530);
  not NOT_12511(g29631,II39011);
  not NOT_12512(II39014,g29535);
  not NOT_12513(g29632,II39014);
  not NOT_12514(II39017,g29542);
  not NOT_12515(g29633,II39017);
  not NOT_12516(II39020,g29499);
  not NOT_12517(g29634,II39020);
  not NOT_12518(II39023,g29508);
  not NOT_12519(g29635,II39023);
  not NOT_12520(II39026,g29510);
  not NOT_12521(g29636,II39026);
  not NOT_12522(II39029,g29512);
  not NOT_12523(g29637,II39029);
  not NOT_12524(II39032,g29537);
  not NOT_12525(g29638,II39032);
  not NOT_12526(II39035,g29544);
  not NOT_12527(g29639,II39035);
  not NOT_12528(II39038,g29551);
  not NOT_12529(g29640,II39038);
  not NOT_12530(II39041,g29501);
  not NOT_12531(g29641,II39041);
  not NOT_12532(II39044,g29511);
  not NOT_12533(g29642,II39044);
  not NOT_12534(II39047,g29513);
  not NOT_12535(g29643,II39047);
  not NOT_12536(II39050,g29515);
  not NOT_12537(g29644,II39050);
  not NOT_12538(II39053,g29546);
  not NOT_12539(g29645,II39053);
  not NOT_12540(II39056,g29554);
  not NOT_12541(g29646,II39056);
  not NOT_12542(II39059,g29561);
  not NOT_12543(g29647,II39059);
  not NOT_12544(II39062,g29504);
  not NOT_12545(g29648,II39062);
  not NOT_12546(II39065,g29514);
  not NOT_12547(g29649,II39065);
  not NOT_12548(II39068,g29516);
  not NOT_12549(g29650,II39068);
  not NOT_12550(II39071,g29517);
  not NOT_12551(g29651,II39071);
  not NOT_12552(II39074,g29556);
  not NOT_12553(g29652,II39074);
  not NOT_12554(II39077,g29563);
  not NOT_12555(g29653,II39077);
  not NOT_12556(II39080,g29568);
  not NOT_12557(g29654,II39080);
  not NOT_12558(II39083,g29519);
  not NOT_12559(g29655,II39083);
  not NOT_12560(II39086,g29497);
  not NOT_12561(g29656,II39086);
  not NOT_12562(II39089,g29495);
  not NOT_12563(g29657,II39089);
  not NOT_12564(g29658,g29574);
  not NOT_12565(g29659,g29571);
  not NOT_12566(g29660,g29578);
  not NOT_12567(g29661,g29576);
  not NOT_12568(g29662,g29570);
  not NOT_12569(g29664,g29552);
  not NOT_12570(g29666,g29577);
  not NOT_12571(g29668,g29569);
  not NOT_12572(g29673,g29583);
  not NOT_12573(II39121,g29579);
  not NOT_12574(g29689,II39121);
  not NOT_12575(II39124,g29606);
  not NOT_12576(g29690,II39124);
  not NOT_12577(II39127,g29608);
  not NOT_12578(g29691,II39127);
  not NOT_12579(II39130,g29580);
  not NOT_12580(g29692,II39130);
  not NOT_12581(II39133,g29609);
  not NOT_12582(g29693,II39133);
  not NOT_12583(II39136,g29611);
  not NOT_12584(g29694,II39136);
  not NOT_12585(II39139,g29612);
  not NOT_12586(g29695,II39139);
  not NOT_12587(II39142,g29581);
  not NOT_12588(g29696,II39142);
  not NOT_12589(II39145,g29613);
  not NOT_12590(g29697,II39145);
  not NOT_12591(II39148,g29616);
  not NOT_12592(g29698,II39148);
  not NOT_12593(II39151,g29617);
  not NOT_12594(g29699,II39151);
  not NOT_12595(II39154,g29582);
  not NOT_12596(g29700,II39154);
  not NOT_12597(II39157,g29618);
  not NOT_12598(g29701,II39157);
  not NOT_12599(II39160,g29620);
  not NOT_12600(g29702,II39160);
  not NOT_12601(II39164,g29621);
  not NOT_12602(g29704,II39164);
  not NOT_12603(II39168,g29623);
  not NOT_12604(g29708,II39168);
  not NOT_12605(g29716,g29498);
  not NOT_12606(g29724,g29500);
  not NOT_12607(g29726,g29503);
  not NOT_12608(g29739,g29505);
  not NOT_12609(II39234,g29689);
  not NOT_12610(g29794,II39234);
  not NOT_12611(II39237,g29690);
  not NOT_12612(g29795,II39237);
  not NOT_12613(II39240,g29691);
  not NOT_12614(g29796,II39240);
  not NOT_12615(II39243,g29694);
  not NOT_12616(g29797,II39243);
  not NOT_12617(II39246,g29692);
  not NOT_12618(g29798,II39246);
  not NOT_12619(II39249,g29693);
  not NOT_12620(g29799,II39249);
  not NOT_12621(II39252,g29695);
  not NOT_12622(g29800,II39252);
  not NOT_12623(II39255,g29698);
  not NOT_12624(g29801,II39255);
  not NOT_12625(II39258,g29696);
  not NOT_12626(g29802,II39258);
  not NOT_12627(II39261,g29697);
  not NOT_12628(g29803,II39261);
  not NOT_12629(II39264,g29699);
  not NOT_12630(g29804,II39264);
  not NOT_12631(II39267,g29702);
  not NOT_12632(g29805,II39267);
  not NOT_12633(II39270,g29700);
  not NOT_12634(g29806,II39270);
  not NOT_12635(II39273,g29701);
  not NOT_12636(g29807,II39273);
  not NOT_12637(II39276,g29704);
  not NOT_12638(g29808,II39276);
  not NOT_12639(II39279,g29708);
  not NOT_12640(g29809,II39279);
  not NOT_12641(g29823,g29663);
  not NOT_12642(g29829,g29665);
  not NOT_12643(g29835,g29667);
  not NOT_12644(g29840,g29669);
  not NOT_12645(g29844,g29670);
  not NOT_12646(g29848,g29761);
  not NOT_12647(g29849,g29671);
  not NOT_12648(g29853,g29672);
  not NOT_12649(g29857,g29676);
  not NOT_12650(g29861,g29677);
  not NOT_12651(g29865,g29678);
  not NOT_12652(g29869,g29679);
  not NOT_12653(g29873,g29680);
  not NOT_12654(g29877,g29681);
  not NOT_12655(g29881,g29682);
  not NOT_12656(g29885,g29683);
  not NOT_12657(g29889,g29684);
  not NOT_12658(g29893,g29685);
  not NOT_12659(g29897,g29686);
  not NOT_12660(g29901,g29687);
  not NOT_12661(g29905,g29688);
  not NOT_12662(II39398,g29664);
  not NOT_12663(g29932,II39398);
  not NOT_12664(II39401,g29662);
  not NOT_12665(g29933,II39401);
  not NOT_12666(II39404,g29661);
  not NOT_12667(g29934,II39404);
  not NOT_12668(II39407,g29660);
  not NOT_12669(g29935,II39407);
  not NOT_12670(II39411,g29659);
  not NOT_12671(g29937,II39411);
  not NOT_12672(II39414,g29658);
  not NOT_12673(g29938,II39414);
  not NOT_12674(II39418,g29668);
  not NOT_12675(g29940,II39418);
  not NOT_12676(II39423,g29666);
  not NOT_12677(g29943,II39423);
  not NOT_12678(II39454,g29940);
  not NOT_12679(g29972,II39454);
  not NOT_12680(II39457,g29943);
  not NOT_12681(g29973,II39457);
  not NOT_12682(II39460,g29932);
  not NOT_12683(g29974,II39460);
  not NOT_12684(II39463,g29933);
  not NOT_12685(g29975,II39463);
  not NOT_12686(II39466,g29934);
  not NOT_12687(g29976,II39466);
  not NOT_12688(II39469,g29935);
  not NOT_12689(g29977,II39469);
  not NOT_12690(II39472,g29937);
  not NOT_12691(g29978,II39472);
  not NOT_12692(II39475,g29938);
  not NOT_12693(g29979,II39475);
  not NOT_12694(g30036,g29912);
  not NOT_12695(g30040,g29914);
  not NOT_12696(g30044,g29916);
  not NOT_12697(g30048,g29920);
  not NOT_12698(II39550,g29848);
  not NOT_12699(g30052,II39550);
  not NOT_12700(II39573,g29936);
  not NOT_12701(g30076,II39573);
  not NOT_12702(II39577,g29939);
  not NOT_12703(g30078,II39577);
  not NOT_12704(II39585,g29941);
  not NOT_12705(g30084,II39585);
  not NOT_12706(II39622,g30052);
  not NOT_12707(g30119,II39622);
  not NOT_12708(II39625,g30076);
  not NOT_12709(g30120,II39625);
  not NOT_12710(II39628,g30078);
  not NOT_12711(g30121,II39628);
  not NOT_12712(II39631,g30084);
  not NOT_12713(g30122,II39631);
  not NOT_12714(II39635,g30055);
  not NOT_12715(g30124,II39635);
  not NOT_12716(II39638,g30056);
  not NOT_12717(g30125,II39638);
  not NOT_12718(II39641,g30057);
  not NOT_12719(g30126,II39641);
  not NOT_12720(II39647,g30058);
  not NOT_12721(g30130,II39647);
  not NOT_12722(g30134,g30010);
  not NOT_12723(g30139,g30011);
  not NOT_12724(g30143,g30012);
  not NOT_12725(g30147,g30013);
  not NOT_12726(g30151,g30014);
  not NOT_12727(g30155,g30015);
  not NOT_12728(g30159,g30016);
  not NOT_12729(g30163,g30017);
  not NOT_12730(g30167,g30018);
  not NOT_12731(g30171,g30019);
  not NOT_12732(g30175,g30020);
  not NOT_12733(g30179,g30021);
  not NOT_12734(g30183,g30022);
  not NOT_12735(g30187,g30023);
  not NOT_12736(g30191,g30024);
  not NOT_12737(g30195,g30025);
  not NOT_12738(g30199,g30026);
  not NOT_12739(g30203,g30027);
  not NOT_12740(g30207,g30028);
  not NOT_12741(g30211,g30029);
  not NOT_12742(II39674,g30072);
  not NOT_12743(g30215,II39674);
  not NOT_12744(g30229,g30030);
  not NOT_12745(g30233,g30031);
  not NOT_12746(g30237,g30032);
  not NOT_12747(g30241,g30033);
  not NOT_12748(II39761,g30072);
  not NOT_12749(g30306,II39761);
  not NOT_12750(II39764,g30060);
  not NOT_12751(g30307,II39764);
  not NOT_12752(II39767,g30061);
  not NOT_12753(g30308,II39767);
  not NOT_12754(II39770,g30063);
  not NOT_12755(g30309,II39770);
  not NOT_12756(II39773,g30064);
  not NOT_12757(g30310,II39773);
  not NOT_12758(II39776,g30066);
  not NOT_12759(g30311,II39776);
  not NOT_12760(II39779,g30053);
  not NOT_12761(g30312,II39779);
  not NOT_12762(II39782,g30054);
  not NOT_12763(g30313,II39782);
  not NOT_12764(II39785,g30124);
  not NOT_12765(g30314,II39785);
  not NOT_12766(II39788,g30125);
  not NOT_12767(g30315,II39788);
  not NOT_12768(II39791,g30126);
  not NOT_12769(g30316,II39791);
  not NOT_12770(II39794,g30130);
  not NOT_12771(g30317,II39794);
  not NOT_12772(II39797,g30307);
  not NOT_12773(g30318,II39797);
  not NOT_12774(II39800,g30309);
  not NOT_12775(g30319,II39800);
  not NOT_12776(II39803,g30308);
  not NOT_12777(g30320,II39803);
  not NOT_12778(II39806,g30310);
  not NOT_12779(g30321,II39806);
  not NOT_12780(II39809,g30311);
  not NOT_12781(g30322,II39809);
  not NOT_12782(II39812,g30312);
  not NOT_12783(g30323,II39812);
  not NOT_12784(II39815,g30313);
  not NOT_12785(g30324,II39815);
  not NOT_12786(II39818,g30215);
  not NOT_12787(g30325,II39818);
  not NOT_12788(II39821,g30267);
  not NOT_12789(g30326,II39821);
  not NOT_12790(II39825,g30268);
  not NOT_12791(g30328,II39825);
  not NOT_12792(II39828,g30269);
  not NOT_12793(g30329,II39828);
  not NOT_12794(II39832,g30270);
  not NOT_12795(g30331,II39832);
  not NOT_12796(II39835,g30271);
  not NOT_12797(g30332,II39835);
  not NOT_12798(II39840,g30272);
  not NOT_12799(g30335,II39840);
  not NOT_12800(II39843,g30273);
  not NOT_12801(g30336,II39843);
  not NOT_12802(II39848,g30274);
  not NOT_12803(g30339,II39848);
  not NOT_12804(II39853,g30275);
  not NOT_12805(g30342,II39853);
  not NOT_12806(II39856,g30276);
  not NOT_12807(g30343,II39856);
  not NOT_12808(II39859,g30277);
  not NOT_12809(g30344,II39859);
  not NOT_12810(II39863,g30278);
  not NOT_12811(g30346,II39863);
  not NOT_12812(II39866,g30279);
  not NOT_12813(g30347,II39866);
  not NOT_12814(II39870,g30280);
  not NOT_12815(g30349,II39870);
  not NOT_12816(II39873,g30281);
  not NOT_12817(g30350,II39873);
  not NOT_12818(II39878,g30282);
  not NOT_12819(g30353,II39878);
  not NOT_12820(II39881,g30283);
  not NOT_12821(g30354,II39881);
  not NOT_12822(II39886,g30284);
  not NOT_12823(g30357,II39886);
  not NOT_12824(II39889,g30285);
  not NOT_12825(g30358,II39889);
  not NOT_12826(II39892,g30286);
  not NOT_12827(g30359,II39892);
  not NOT_12828(II39895,g30287);
  not NOT_12829(g30360,II39895);
  not NOT_12830(II39899,g30288);
  not NOT_12831(g30362,II39899);
  not NOT_12832(II39902,g30289);
  not NOT_12833(g30363,II39902);
  not NOT_12834(II39906,g30290);
  not NOT_12835(g30365,II39906);
  not NOT_12836(II39909,g30291);
  not NOT_12837(g30366,II39909);
  not NOT_12838(II39913,g30292);
  not NOT_12839(g30368,II39913);
  not NOT_12840(II39916,g30293);
  not NOT_12841(g30369,II39916);
  not NOT_12842(II39919,g30294);
  not NOT_12843(g30370,II39919);
  not NOT_12844(II39922,g30295);
  not NOT_12845(g30371,II39922);
  not NOT_12846(II39926,g30296);
  not NOT_12847(g30373,II39926);
  not NOT_12848(II39930,g30297);
  not NOT_12849(g30375,II39930);
  not NOT_12850(II39933,g30298);
  not NOT_12851(g30376,II39933);
  not NOT_12852(II39936,g30299);
  not NOT_12853(g30377,II39936);
  not NOT_12854(II39939,g30300);
  not NOT_12855(g30378,II39939);
  not NOT_12856(II39942,g30301);
  not NOT_12857(g30379,II39942);
  not NOT_12858(II39945,g30302);
  not NOT_12859(g30380,II39945);
  not NOT_12860(II39948,g30303);
  not NOT_12861(g30381,II39948);
  not NOT_12862(II39951,g30304);
  not NOT_12863(g30382,II39951);
  not NOT_12864(g30383,g30306);
  not NOT_12865(II39976,g30245);
  not NOT_12866(g30408,II39976);
  not NOT_12867(II39982,g30305);
  not NOT_12868(g30412,II39982);
  not NOT_12869(II39985,g30246);
  not NOT_12870(g30435,II39985);
  not NOT_12871(II39991,g30247);
  not NOT_12872(g30439,II39991);
  not NOT_12873(II39997,g30248);
  not NOT_12874(g30443,II39997);
  not NOT_12875(II40002,g30249);
  not NOT_12876(g30446,II40002);
  not NOT_12877(II40008,g30250);
  not NOT_12878(g30450,II40008);
  not NOT_12879(II40016,g30251);
  not NOT_12880(g30456,II40016);
  not NOT_12881(II40021,g30252);
  not NOT_12882(g30459,II40021);
  not NOT_12883(II40027,g30253);
  not NOT_12884(g30463,II40027);
  not NOT_12885(II40032,g30254);
  not NOT_12886(g30466,II40032);
  not NOT_12887(II40039,g30255);
  not NOT_12888(g30471,II40039);
  not NOT_12889(II40044,g30256);
  not NOT_12890(g30474,II40044);
  not NOT_12891(II40051,g30257);
  not NOT_12892(g30479,II40051);
  not NOT_12893(II40054,g30258);
  not NOT_12894(g30480,II40054);
  not NOT_12895(II40059,g30259);
  not NOT_12896(g30483,II40059);
  not NOT_12897(II40066,g30260);
  not NOT_12898(g30488,II40066);
  not NOT_12899(II40071,g30261);
  not NOT_12900(g30491,II40071);
  not NOT_12901(II40075,g30262);
  not NOT_12902(g30493,II40075);
  not NOT_12903(II40078,g30263);
  not NOT_12904(g30494,II40078);
  not NOT_12905(II40083,g30264);
  not NOT_12906(g30497,II40083);
  not NOT_12907(II40086,g30265);
  not NOT_12908(g30498,II40086);
  not NOT_12909(II40091,g30266);
  not NOT_12910(g30501,II40091);
  not NOT_12911(II40098,g30491);
  not NOT_12912(g30506,II40098);
  not NOT_12913(II40101,g30326);
  not NOT_12914(g30507,II40101);
  not NOT_12915(II40104,g30342);
  not NOT_12916(g30508,II40104);
  not NOT_12917(II40107,g30343);
  not NOT_12918(g30509,II40107);
  not NOT_12919(II40110,g30357);
  not NOT_12920(g30510,II40110);
  not NOT_12921(II40113,g30368);
  not NOT_12922(g30511,II40113);
  not NOT_12923(II40116,g30408);
  not NOT_12924(g30512,II40116);
  not NOT_12925(II40119,g30435);
  not NOT_12926(g30513,II40119);
  not NOT_12927(II40122,g30443);
  not NOT_12928(g30514,II40122);
  not NOT_12929(II40125,g30466);
  not NOT_12930(g30515,II40125);
  not NOT_12931(II40128,g30479);
  not NOT_12932(g30516,II40128);
  not NOT_12933(II40131,g30493);
  not NOT_12934(g30517,II40131);
  not NOT_12935(II40134,g30480);
  not NOT_12936(g30518,II40134);
  not NOT_12937(II40137,g30494);
  not NOT_12938(g30519,II40137);
  not NOT_12939(II40140,g30328);
  not NOT_12940(g30520,II40140);
  not NOT_12941(II40143,g30329);
  not NOT_12942(g30521,II40143);
  not NOT_12943(II40146,g30344);
  not NOT_12944(g30522,II40146);
  not NOT_12945(II40149,g30358);
  not NOT_12946(g30523,II40149);
  not NOT_12947(II40152,g30359);
  not NOT_12948(g30524,II40152);
  not NOT_12949(II40155,g30369);
  not NOT_12950(g30525,II40155);
  not NOT_12951(II40158,g30376);
  not NOT_12952(g30526,II40158);
  not NOT_12953(II40161,g30439);
  not NOT_12954(g30527,II40161);
  not NOT_12955(II40164,g30446);
  not NOT_12956(g30528,II40164);
  not NOT_12957(II40167,g30456);
  not NOT_12958(g30529,II40167);
  not NOT_12959(II40170,g30483);
  not NOT_12960(g30530,II40170);
  not NOT_12961(II40173,g30497);
  not NOT_12962(g30531,II40173);
  not NOT_12963(II40176,g30331);
  not NOT_12964(g30532,II40176);
  not NOT_12965(II40179,g30498);
  not NOT_12966(g30533,II40179);
  not NOT_12967(II40182,g30332);
  not NOT_12968(g30534,II40182);
  not NOT_12969(II40185,g30346);
  not NOT_12970(g30535,II40185);
  not NOT_12971(II40188,g30347);
  not NOT_12972(g30536,II40188);
  not NOT_12973(II40191,g30360);
  not NOT_12974(g30537,II40191);
  not NOT_12975(II40194,g30370);
  not NOT_12976(g30538,II40194);
  not NOT_12977(II40197,g30371);
  not NOT_12978(g30539,II40197);
  not NOT_12979(II40200,g30377);
  not NOT_12980(g30540,II40200);
  not NOT_12981(II40203,g30380);
  not NOT_12982(g30541,II40203);
  not NOT_12983(II40206,g30450);
  not NOT_12984(g30542,II40206);
  not NOT_12985(II40209,g30459);
  not NOT_12986(g30543,II40209);
  not NOT_12987(II40212,g30471);
  not NOT_12988(g30544,II40212);
  not NOT_12989(II40215,g30501);
  not NOT_12990(g30545,II40215);
  not NOT_12991(II40218,g30335);
  not NOT_12992(g30546,II40218);
  not NOT_12993(II40221,g30349);
  not NOT_12994(g30547,II40221);
  not NOT_12995(II40224,g30336);
  not NOT_12996(g30548,II40224);
  not NOT_12997(II40227,g30350);
  not NOT_12998(g30549,II40227);
  not NOT_12999(II40230,g30362);
  not NOT_13000(g30550,II40230);
  not NOT_13001(II40233,g30363);
  not NOT_13002(g30551,II40233);
  not NOT_13003(II40236,g30373);
  not NOT_13004(g30552,II40236);
  not NOT_13005(II40239,g30378);
  not NOT_13006(g30553,II40239);
  not NOT_13007(II40242,g30379);
  not NOT_13008(g30554,II40242);
  not NOT_13009(II40245,g30381);
  not NOT_13010(g30555,II40245);
  not NOT_13011(II40248,g30382);
  not NOT_13012(g30556,II40248);
  not NOT_13013(II40251,g30463);
  not NOT_13014(g30557,II40251);
  not NOT_13015(II40254,g30474);
  not NOT_13016(g30558,II40254);
  not NOT_13017(II40257,g30488);
  not NOT_13018(g30559,II40257);
  not NOT_13019(II40260,g30339);
  not NOT_13020(g30560,II40260);
  not NOT_13021(II40263,g30353);
  not NOT_13022(g30561,II40263);
  not NOT_13023(II40266,g30365);
  not NOT_13024(g30562,II40266);
  not NOT_13025(II40269,g30354);
  not NOT_13026(g30563,II40269);
  not NOT_13027(II40272,g30366);
  not NOT_13028(g30564,II40272);
  not NOT_13029(II40275,g30375);
  not NOT_13030(g30565,II40275);
  not NOT_13031(g30567,g30403);
  not NOT_13032(g30568,g30402);
  not NOT_13033(g30569,g30406);
  not NOT_13034(g30570,g30404);
  not NOT_13035(g30571,g30401);
  not NOT_13036(g30572,g30399);
  not NOT_13037(g30573,g30405);
  not NOT_13038(g30574,g30400);
  not NOT_13039(g30575,g30412);
  not NOT_13040(II40288,g30455);
  not NOT_13041(g30578,II40288);
  not NOT_13042(II40291,g30468);
  not NOT_13043(g30579,II40291);
  not NOT_13044(II40294,g30470);
  not NOT_13045(g30580,II40294);
  not NOT_13046(II40297,g30482);
  not NOT_13047(g30581,II40297);
  not NOT_13048(II40300,g30485);
  not NOT_13049(g30582,II40300);
  not NOT_13050(II40303,g30487);
  not NOT_13051(g30583,II40303);
  not NOT_13052(II40307,g30500);
  not NOT_13053(g30585,II40307);
  not NOT_13054(II40310,g30503);
  not NOT_13055(g30586,II40310);
  not NOT_13056(II40313,g30505);
  not NOT_13057(g30587,II40313);
  not NOT_13058(II40317,g30338);
  not NOT_13059(g30591,II40317);
  not NOT_13060(II40320,g30341);
  not NOT_13061(g30592,II40320);
  not NOT_13062(II40326,g30356);
  not NOT_13063(g30600,II40326);
  not NOT_13064(II40420,g30578);
  not NOT_13065(g30710,II40420);
  not NOT_13066(II40423,g30579);
  not NOT_13067(g30711,II40423);
  not NOT_13068(II40426,g30581);
  not NOT_13069(g30712,II40426);
  not NOT_13070(II40429,g30580);
  not NOT_13071(g30713,II40429);
  not NOT_13072(II40432,g30582);
  not NOT_13073(g30714,II40432);
  not NOT_13074(II40435,g30585);
  not NOT_13075(g30715,II40435);
  not NOT_13076(II40438,g30583);
  not NOT_13077(g30716,II40438);
  not NOT_13078(II40441,g30586);
  not NOT_13079(g30717,II40441);
  not NOT_13080(II40444,g30591);
  not NOT_13081(g30718,II40444);
  not NOT_13082(II40447,g30587);
  not NOT_13083(g30719,II40447);
  not NOT_13084(II40450,g30592);
  not NOT_13085(g30720,II40450);
  not NOT_13086(II40453,g30600);
  not NOT_13087(g30721,II40453);
  not NOT_13088(II40456,g30668);
  not NOT_13089(g30722,II40456);
  not NOT_13090(II40459,g30669);
  not NOT_13091(g30723,II40459);
  not NOT_13092(II40462,g30670);
  not NOT_13093(g30724,II40462);
  not NOT_13094(II40465,g30671);
  not NOT_13095(g30725,II40465);
  not NOT_13096(II40468,g30672);
  not NOT_13097(g30726,II40468);
  not NOT_13098(II40471,g30673);
  not NOT_13099(g30727,II40471);
  not NOT_13100(II40475,g30674);
  not NOT_13101(g30729,II40475);
  not NOT_13102(II40478,g30675);
  not NOT_13103(g30730,II40478);
  not NOT_13104(II40481,g30676);
  not NOT_13105(g30731,II40481);
  not NOT_13106(II40484,g30677);
  not NOT_13107(g30732,II40484);
  not NOT_13108(II40487,g30678);
  not NOT_13109(g30733,II40487);
  not NOT_13110(II40490,g30679);
  not NOT_13111(g30734,II40490);
  not NOT_13112(II40495,g30680);
  not NOT_13113(g30737,II40495);
  not NOT_13114(II40498,g30681);
  not NOT_13115(g30738,II40498);
  not NOT_13116(II40501,g30682);
  not NOT_13117(g30739,II40501);
  not NOT_13118(II40504,g30683);
  not NOT_13119(g30740,II40504);
  not NOT_13120(II40507,g30684);
  not NOT_13121(g30741,II40507);
  not NOT_13122(II40510,g30686);
  not NOT_13123(g30742,II40510);
  not NOT_13124(II40515,g30687);
  not NOT_13125(g30745,II40515);
  not NOT_13126(II40518,g30688);
  not NOT_13127(g30746,II40518);
  not NOT_13128(II40521,g30689);
  not NOT_13129(g30747,II40521);
  not NOT_13130(II40524,g30690);
  not NOT_13131(g30748,II40524);
  not NOT_13132(II40527,g30691);
  not NOT_13133(g30749,II40527);
  not NOT_13134(II40531,g30692);
  not NOT_13135(g30751,II40531);
  not NOT_13136(II40534,g30693);
  not NOT_13137(g30752,II40534);
  not NOT_13138(II40537,g30694);
  not NOT_13139(g30753,II40537);
  not NOT_13140(II40542,g30695);
  not NOT_13141(g30756,II40542);
  not NOT_13142(g30765,g30685);
  not NOT_13143(II40555,g30699);
  not NOT_13144(g30767,II40555);
  not NOT_13145(II40565,g30700);
  not NOT_13146(g30769,II40565);
  not NOT_13147(II40568,g30701);
  not NOT_13148(g30770,II40568);
  not NOT_13149(II40578,g30702);
  not NOT_13150(g30772,II40578);
  not NOT_13151(II40581,g30703);
  not NOT_13152(g30773,II40581);
  not NOT_13153(II40584,g30704);
  not NOT_13154(g30774,II40584);
  not NOT_13155(II40594,g30705);
  not NOT_13156(g30776,II40594);
  not NOT_13157(II40597,g30706);
  not NOT_13158(g30777,II40597);
  not NOT_13159(II40600,g30707);
  not NOT_13160(g30778,II40600);
  not NOT_13161(II40611,g30708);
  not NOT_13162(g30781,II40611);
  not NOT_13163(II40614,g30709);
  not NOT_13164(g30782,II40614);
  not NOT_13165(II40618,g30566);
  not NOT_13166(g30784,II40618);
  not NOT_13167(II40634,g30571);
  not NOT_13168(g30792,II40634);
  not NOT_13169(II40637,g30570);
  not NOT_13170(g30793,II40637);
  not NOT_13171(II40640,g30569);
  not NOT_13172(g30794,II40640);
  not NOT_13173(II40643,g30568);
  not NOT_13174(g30795,II40643);
  not NOT_13175(II40647,g30567);
  not NOT_13176(g30797,II40647);
  not NOT_13177(II40651,g30574);
  not NOT_13178(g30799,II40651);
  not NOT_13179(II40654,g30573);
  not NOT_13180(g30800,II40654);
  not NOT_13181(II40658,g30572);
  not NOT_13182(g30802,II40658);
  not NOT_13183(II40661,g30635);
  not NOT_13184(g30803,II40661);
  not NOT_13185(II40664,g30636);
  not NOT_13186(g30804,II40664);
  not NOT_13187(II40667,g30637);
  not NOT_13188(g30805,II40667);
  not NOT_13189(II40670,g30638);
  not NOT_13190(g30806,II40670);
  not NOT_13191(II40673,g30639);
  not NOT_13192(g30807,II40673);
  not NOT_13193(II40676,g30640);
  not NOT_13194(g30808,II40676);
  not NOT_13195(II40679,g30641);
  not NOT_13196(g30809,II40679);
  not NOT_13197(II40682,g30642);
  not NOT_13198(g30810,II40682);
  not NOT_13199(II40685,g30643);
  not NOT_13200(g30811,II40685);
  not NOT_13201(II40688,g30644);
  not NOT_13202(g30812,II40688);
  not NOT_13203(II40691,g30645);
  not NOT_13204(g30813,II40691);
  not NOT_13205(II40694,g30646);
  not NOT_13206(g30814,II40694);
  not NOT_13207(II40697,g30647);
  not NOT_13208(g30815,II40697);
  not NOT_13209(II40700,g30648);
  not NOT_13210(g30816,II40700);
  not NOT_13211(II40703,g30649);
  not NOT_13212(g30817,II40703);
  not NOT_13213(II40706,g30650);
  not NOT_13214(g30818,II40706);
  not NOT_13215(II40709,g30651);
  not NOT_13216(g30819,II40709);
  not NOT_13217(II40712,g30652);
  not NOT_13218(g30820,II40712);
  not NOT_13219(II40715,g30653);
  not NOT_13220(g30821,II40715);
  not NOT_13221(II40718,g30654);
  not NOT_13222(g30822,II40718);
  not NOT_13223(II40721,g30655);
  not NOT_13224(g30823,II40721);
  not NOT_13225(II40724,g30656);
  not NOT_13226(g30824,II40724);
  not NOT_13227(II40727,g30657);
  not NOT_13228(g30825,II40727);
  not NOT_13229(II40730,g30658);
  not NOT_13230(g30826,II40730);
  not NOT_13231(II40733,g30659);
  not NOT_13232(g30827,II40733);
  not NOT_13233(II40736,g30660);
  not NOT_13234(g30828,II40736);
  not NOT_13235(II40739,g30661);
  not NOT_13236(g30829,II40739);
  not NOT_13237(II40742,g30662);
  not NOT_13238(g30830,II40742);
  not NOT_13239(II40745,g30663);
  not NOT_13240(g30831,II40745);
  not NOT_13241(II40748,g30664);
  not NOT_13242(g30832,II40748);
  not NOT_13243(II40751,g30665);
  not NOT_13244(g30833,II40751);
  not NOT_13245(II40754,g30666);
  not NOT_13246(g30834,II40754);
  not NOT_13247(II40757,g30667);
  not NOT_13248(g30835,II40757);
  not NOT_13249(II40760,g30722);
  not NOT_13250(g30836,II40760);
  not NOT_13251(II40763,g30729);
  not NOT_13252(g30837,II40763);
  not NOT_13253(II40766,g30737);
  not NOT_13254(g30838,II40766);
  not NOT_13255(II40769,g30803);
  not NOT_13256(g30839,II40769);
  not NOT_13257(II40772,g30804);
  not NOT_13258(g30840,II40772);
  not NOT_13259(II40775,g30807);
  not NOT_13260(g30841,II40775);
  not NOT_13261(II40778,g30805);
  not NOT_13262(g30842,II40778);
  not NOT_13263(II40781,g30808);
  not NOT_13264(g30843,II40781);
  not NOT_13265(II40784,g30813);
  not NOT_13266(g30844,II40784);
  not NOT_13267(II40787,g30809);
  not NOT_13268(g30845,II40787);
  not NOT_13269(II40790,g30814);
  not NOT_13270(g30846,II40790);
  not NOT_13271(II40793,g30821);
  not NOT_13272(g30847,II40793);
  not NOT_13273(II40796,g30829);
  not NOT_13274(g30848,II40796);
  not NOT_13275(II40799,g30723);
  not NOT_13276(g30849,II40799);
  not NOT_13277(II40802,g30730);
  not NOT_13278(g30850,II40802);
  not NOT_13279(II40805,g30767);
  not NOT_13280(g30851,II40805);
  not NOT_13281(II40808,g30769);
  not NOT_13282(g30852,II40808);
  not NOT_13283(II40811,g30772);
  not NOT_13284(g30853,II40811);
  not NOT_13285(II40814,g30731);
  not NOT_13286(g30854,II40814);
  not NOT_13287(II40817,g30738);
  not NOT_13288(g30855,II40817);
  not NOT_13289(II40820,g30745);
  not NOT_13290(g30856,II40820);
  not NOT_13291(II40823,g30806);
  not NOT_13292(g30857,II40823);
  not NOT_13293(II40826,g30810);
  not NOT_13294(g30858,II40826);
  not NOT_13295(II40829,g30815);
  not NOT_13296(g30859,II40829);
  not NOT_13297(II40832,g30811);
  not NOT_13298(g30860,II40832);
  not NOT_13299(II40835,g30816);
  not NOT_13300(g30861,II40835);
  not NOT_13301(II40838,g30822);
  not NOT_13302(g30862,II40838);
  not NOT_13303(II40841,g30817);
  not NOT_13304(g30863,II40841);
  not NOT_13305(II40844,g30823);
  not NOT_13306(g30864,II40844);
  not NOT_13307(II40847,g30830);
  not NOT_13308(g30865,II40847);
  not NOT_13309(II40850,g30724);
  not NOT_13310(g30866,II40850);
  not NOT_13311(II40853,g30732);
  not NOT_13312(g30867,II40853);
  not NOT_13313(II40856,g30739);
  not NOT_13314(g30868,II40856);
  not NOT_13315(II40859,g30770);
  not NOT_13316(g30869,II40859);
  not NOT_13317(II40862,g30773);
  not NOT_13318(g30870,II40862);
  not NOT_13319(II40865,g30776);
  not NOT_13320(g30871,II40865);
  not NOT_13321(II40868,g30740);
  not NOT_13322(g30872,II40868);
  not NOT_13323(II40871,g30746);
  not NOT_13324(g30873,II40871);
  not NOT_13325(II40874,g30751);
  not NOT_13326(g30874,II40874);
  not NOT_13327(II40877,g30812);
  not NOT_13328(g30875,II40877);
  not NOT_13329(II40880,g30818);
  not NOT_13330(g30876,II40880);
  not NOT_13331(II40883,g30824);
  not NOT_13332(g30877,II40883);
  not NOT_13333(II40886,g30819);
  not NOT_13334(g30878,II40886);
  not NOT_13335(II40889,g30825);
  not NOT_13336(g30879,II40889);
  not NOT_13337(II40892,g30831);
  not NOT_13338(g30880,II40892);
  not NOT_13339(II40895,g30826);
  not NOT_13340(g30881,II40895);
  not NOT_13341(II40898,g30832);
  not NOT_13342(g30882,II40898);
  not NOT_13343(II40901,g30725);
  not NOT_13344(g30883,II40901);
  not NOT_13345(II40904,g30733);
  not NOT_13346(g30884,II40904);
  not NOT_13347(II40907,g30741);
  not NOT_13348(g30885,II40907);
  not NOT_13349(II40910,g30747);
  not NOT_13350(g30886,II40910);
  not NOT_13351(II40913,g30774);
  not NOT_13352(g30887,II40913);
  not NOT_13353(II40916,g30777);
  not NOT_13354(g30888,II40916);
  not NOT_13355(II40919,g30781);
  not NOT_13356(g30889,II40919);
  not NOT_13357(II40922,g30748);
  not NOT_13358(g30890,II40922);
  not NOT_13359(II40925,g30752);
  not NOT_13360(g30891,II40925);
  not NOT_13361(II40928,g30756);
  not NOT_13362(g30892,II40928);
  not NOT_13363(II40931,g30820);
  not NOT_13364(g30893,II40931);
  not NOT_13365(II40934,g30827);
  not NOT_13366(g30894,II40934);
  not NOT_13367(II40937,g30833);
  not NOT_13368(g30895,II40937);
  not NOT_13369(II40940,g30828);
  not NOT_13370(g30896,II40940);
  not NOT_13371(II40943,g30834);
  not NOT_13372(g30897,II40943);
  not NOT_13373(II40946,g30726);
  not NOT_13374(g30898,II40946);
  not NOT_13375(II40949,g30835);
  not NOT_13376(g30899,II40949);
  not NOT_13377(II40952,g30727);
  not NOT_13378(g30900,II40952);
  not NOT_13379(II40955,g30734);
  not NOT_13380(g30901,II40955);
  not NOT_13381(II40958,g30742);
  not NOT_13382(g30902,II40958);
  not NOT_13383(II40961,g30749);
  not NOT_13384(g30903,II40961);
  not NOT_13385(II40964,g30753);
  not NOT_13386(g30904,II40964);
  not NOT_13387(II40967,g30778);
  not NOT_13388(g30905,II40967);
  not NOT_13389(II40970,g30782);
  not NOT_13390(g30906,II40970);
  not NOT_13391(II40973,g30784);
  not NOT_13392(g30907,II40973);
  not NOT_13393(II40976,g30799);
  not NOT_13394(g30908,II40976);
  not NOT_13395(II40979,g30800);
  not NOT_13396(g30909,II40979);
  not NOT_13397(II40982,g30802);
  not NOT_13398(g30910,II40982);
  not NOT_13399(II40985,g30792);
  not NOT_13400(g30911,II40985);
  not NOT_13401(II40988,g30793);
  not NOT_13402(g30912,II40988);
  not NOT_13403(II40991,g30794);
  not NOT_13404(g30913,II40991);
  not NOT_13405(II40994,g30795);
  not NOT_13406(g30914,II40994);
  not NOT_13407(II40997,g30797);
  not NOT_13408(g30915,II40997);
  not NOT_13409(II41024,g30765);
  not NOT_13410(g30928,II41024);
  not NOT_13411(II41035,g30796);
  not NOT_13412(g30937,II41035);
  not NOT_13413(II41038,g30798);
  not NOT_13414(g30938,II41038);
  not NOT_13415(II41041,g30801);
  not NOT_13416(g30939,II41041);
  not NOT_13417(II41044,g30928);
  not NOT_13418(g30940,II41044);
  not NOT_13419(II41047,g30937);
  not NOT_13420(g30941,II41047);
  not NOT_13421(II41050,g30938);
  not NOT_13422(g30942,II41050);
  not NOT_13423(II41053,g30939);
  not NOT_13424(g30943,II41053);
  not NOT_13425(g30962,g30958);
  not NOT_13426(g30963,g30957);
  not NOT_13427(g30964,g30961);
  not NOT_13428(g30965,g30959);
  not NOT_13429(g30966,g30956);
  not NOT_13430(g30967,g30954);
  not NOT_13431(g30968,g30960);
  not NOT_13432(g30969,g30955);
  not NOT_13433(g30971,g30970);
  not NOT_13434(II41090,g30965);
  not NOT_13435(g30972,II41090);
  not NOT_13436(II41093,g30964);
  not NOT_13437(g30973,II41093);
  not NOT_13438(II41096,g30963);
  not NOT_13439(g30974,II41096);
  not NOT_13440(II41099,g30962);
  not NOT_13441(g30975,II41099);
  not NOT_13442(II41102,g30969);
  not NOT_13443(g30976,II41102);
  not NOT_13444(II41105,g30968);
  not NOT_13445(g30977,II41105);
  not NOT_13446(II41108,g30967);
  not NOT_13447(g30978,II41108);
  not NOT_13448(II41111,g30966);
  not NOT_13449(g30979,II41111);
  not NOT_13450(II41114,g30976);
  not NOT_13451(g30980,II41114);
  not NOT_13452(II41117,g30977);
  not NOT_13453(g30981,II41117);
  not NOT_13454(II41120,g30978);
  not NOT_13455(g30982,II41120);
  not NOT_13456(II41123,g30979);
  not NOT_13457(g30983,II41123);
  not NOT_13458(II41126,g30972);
  not NOT_13459(g30984,II41126);
  not NOT_13460(II41129,g30973);
  not NOT_13461(g30985,II41129);
  not NOT_13462(II41132,g30974);
  not NOT_13463(g30986,II41132);
  not NOT_13464(II41135,g30975);
  not NOT_13465(g30987,II41135);
  not NOT_13466(II41138,g30971);
  not NOT_13467(g30988,II41138);
  not NOT_13468(II41141,g30988);
  not NOT_13469(g30989,II41141);
  and AND2_0(g5630,g325,g349);
  and AND2_1(g5649,g331,g351);
  and AND2_2(g5650,g325,g364);
  and AND2_3(g5658,g1012,g1036);
  and AND2_4(g5676,g337,g353);
  and AND2_5(g5677,g331,g366);
  and AND2_6(g5678,g325,g379);
  and AND2_7(g5687,g1018,g1038);
  and AND2_8(g5688,g1012,g1051);
  and AND2_9(g5696,g1706,g1730);
  and AND2_10(g5709,g337,g368);
  and AND2_11(g5710,g331,g381);
  and AND2_12(g5711,g325,g394);
  and AND2_13(g5728,g1024,g1040);
  and AND2_14(g5729,g1018,g1053);
  and AND2_15(g5730,g1012,g1066);
  and AND2_16(g5739,g1712,g1732);
  and AND2_17(g5740,g1706,g1745);
  and AND2_18(g5748,g2400,g2424);
  and AND2_19(g5757,g337,g383);
  and AND2_20(g5758,g331,g396);
  and AND2_21(g5767,g1024,g1055);
  and AND2_22(g5768,g1018,g1068);
  and AND2_23(g5769,g1012,g1081);
  and AND2_24(g5786,g1718,g1734);
  and AND2_25(g5787,g1712,g1747);
  and AND2_26(g5788,g1706,g1760);
  and AND2_27(g5797,g2406,g2426);
  and AND2_28(g5798,g2400,g2439);
  and AND2_29(g5807,g337,g324);
  and AND2_30(g5816,g1024,g1070);
  and AND2_31(g5817,g1018,g1083);
  and AND2_32(g5826,g1718,g1749);
  and AND2_33(g5827,g1712,g1762);
  and AND2_34(g5828,g1706,g1775);
  and AND2_35(g5845,g2412,g2428);
  and AND2_36(g5846,g2406,g2441);
  and AND2_37(g5847,g2400,g2454);
  and AND2_38(g5863,g1024,g1011);
  and AND2_39(g5872,g1718,g1764);
  and AND2_40(g5873,g1712,g1777);
  and AND2_41(g5882,g2412,g2443);
  and AND2_42(g5883,g2406,g2456);
  and AND2_43(g5884,g2400,g2469);
  and AND2_44(g5910,g1718,g1705);
  and AND2_45(g5919,g2412,g2458);
  and AND2_46(g5920,g2406,g2471);
  and AND2_47(g5949,g2412,g2399);
  and AND2_48(g8327,g3254,g219);
  and AND2_49(g8328,g6314,g225);
  and AND2_50(g8329,g6232,g231);
  and AND2_51(g8339,g6519,g903);
  and AND2_52(g8340,g6369,g909);
  and AND2_53(g8350,g6574,g1594);
  and AND2_54(g8385,g3254,g228);
  and AND2_55(g8386,g6314,g234);
  and AND2_56(g8387,g6232,g240);
  and AND2_57(g8394,g3410,g906);
  and AND2_58(g8395,g6519,g912);
  and AND2_59(g8396,g6369,g918);
  and AND2_60(g8406,g6783,g1597);
  and AND2_61(g8407,g6574,g1603);
  and AND2_62(g8417,g6838,g2288);
  and AND2_63(g8431,g3254,g237);
  and AND2_64(g8432,g6314,g243);
  and AND2_65(g8433,g6232,g249);
  and AND2_66(g8437,g3410,g915);
  and AND2_67(g8438,g6519,g921);
  and AND2_68(g8439,g6369,g927);
  and AND2_69(g8446,g3566,g1600);
  and AND2_70(g8447,g6783,g1606);
  and AND2_71(g8448,g6574,g1612);
  and AND2_72(g8458,g7085,g2291);
  and AND2_73(g8459,g6838,g2297);
  and AND2_74(g8463,g3254,g246);
  and AND2_75(g8464,g6314,g252);
  and AND2_76(g8465,g6232,g258);
  and AND2_77(g8466,g3410,g924);
  and AND2_78(g8467,g6519,g930);
  and AND2_79(g8468,g6369,g936);
  and AND2_80(g8472,g3566,g1609);
  and AND2_81(g8473,g6783,g1615);
  and AND2_82(g8474,g6574,g1621);
  and AND2_83(g8481,g3722,g2294);
  and AND2_84(g8482,g7085,g2300);
  and AND2_85(g8483,g6838,g2306);
  and AND2_86(g8484,g6232,g186);
  and AND2_87(g8485,g3254,g255);
  and AND2_88(g8486,g6314,g261);
  and AND2_89(g8487,g6232,g267);
  and AND2_90(g8488,g3410,g933);
  and AND2_91(g8489,g6519,g939);
  and AND2_92(g8490,g6369,g945);
  and AND2_93(g8491,g3566,g1618);
  and AND2_94(g8492,g6783,g1624);
  and AND2_95(g8493,g6574,g1630);
  and AND2_96(g8497,g3722,g2303);
  and AND2_97(g8498,g7085,g2309);
  and AND2_98(g8499,g6838,g2315);
  and AND2_99(g8500,g6314,g189);
  and AND2_100(g8501,g6232,g195);
  and AND2_101(g8502,g3254,g264);
  and AND2_102(g8503,g6314,g270);
  and AND2_103(g8504,g6369,g873);
  and AND2_104(g8505,g3410,g942);
  and AND2_105(g8506,g6519,g948);
  and AND2_106(g8507,g6369,g954);
  and AND2_107(g8508,g3566,g1627);
  and AND2_108(g8509,g6783,g1633);
  and AND2_109(g8510,g6574,g1639);
  and AND2_110(g8511,g3722,g2312);
  and AND2_111(g8512,g7085,g2318);
  and AND2_112(g8513,g6838,g2324);
  and AND2_113(g8515,g3254,g192);
  and AND2_114(g8516,g6314,g198);
  and AND2_115(g8517,g6232,g204);
  and AND2_116(g8518,g3254,g273);
  and AND2_117(g8519,g6519,g876);
  and AND2_118(g8520,g6369,g882);
  and AND2_119(g8521,g3410,g951);
  and AND2_120(g8522,g6519,g957);
  and AND2_121(g8523,g6574,g1567);
  and AND2_122(g8524,g3566,g1636);
  and AND2_123(g8525,g6783,g1642);
  and AND2_124(g8526,g6574,g1648);
  and AND2_125(g8527,g3722,g2321);
  and AND2_126(g8528,g7085,g2327);
  and AND2_127(g8529,g6838,g2333);
  and AND2_128(g8531,g3254,g201);
  and AND2_129(g8532,g6314,g207);
  and AND2_130(g8534,g3410,g879);
  and AND2_131(g8535,g6519,g885);
  and AND2_132(g8536,g6369,g891);
  and AND2_133(g8537,g3410,g960);
  and AND2_134(g8538,g6783,g1570);
  and AND2_135(g8539,g6574,g1576);
  and AND2_136(g8540,g3566,g1645);
  and AND2_137(g8541,g6783,g1651);
  and AND2_138(g8542,g6838,g2261);
  and AND2_139(g8543,g3722,g2330);
  and AND2_140(g8544,g7085,g2336);
  and AND2_141(g8545,g6838,g2342);
  and AND2_142(g8546,g3254,g210);
  and AND2_143(g8548,g3410,g888);
  and AND2_144(g8549,g6519,g894);
  and AND2_145(g8551,g3566,g1573);
  and AND2_146(g8552,g6783,g1579);
  and AND2_147(g8553,g6574,g1585);
  and AND2_148(g8554,g3566,g1654);
  and AND2_149(g8555,g7085,g2264);
  and AND2_150(g8556,g6838,g2270);
  and AND2_151(g8557,g3722,g2339);
  and AND2_152(g8558,g7085,g2345);
  and AND2_153(g8559,g3410,g897);
  and AND2_154(g8561,g3566,g1582);
  and AND2_155(g8562,g6783,g1588);
  and AND2_156(g8564,g3722,g2267);
  and AND2_157(g8565,g7085,g2273);
  and AND2_158(g8566,g6838,g2279);
  and AND2_159(g8567,g3722,g2348);
  and AND2_160(g8570,g3566,g1591);
  and AND2_161(g8572,g3722,g2276);
  and AND2_162(g8573,g7085,g2282);
  and AND2_163(g8576,g3722,g2285);
  and AND2_164(g8601,g6643,g7153);
  and AND2_165(g8612,g3338,g6908);
  and AND2_166(g8613,g6945,g7349);
  and AND2_167(g8621,g6486,g6672);
  and AND2_168(g8625,g3494,g7158);
  and AND2_169(g8626,g7195,g7479);
  and AND2_170(g8631,g6751,g6974);
  and AND2_171(g8635,g3650,g7354);
  and AND2_172(g8636,g7391,g7535);
  and AND2_173(g8650,g7053,g7224);
  and AND2_174(g8654,g3806,g7484);
  and AND2_175(g8666,g7303,g7420);
  and AND2_176(g8676,g6643,g7838);
  and AND2_177(g8687,g3338,g7827);
  and AND2_178(g8688,g6945,g7858);
  and AND2_179(g8703,g6486,g7819);
  and AND2_180(g8704,g6643,g7996);
  and AND2_181(g8705,g3494,g7842);
  and AND2_182(g8706,g7195,g7888);
  and AND2_183(g8717,g3338,g7953);
  and AND2_184(g8722,g6751,g7830);
  and AND2_185(g8723,g6945,g8071);
  and AND2_186(g8724,g3650,g7862);
  and AND2_187(g8725,g7391,g7912);
  and AND2_188(g8751,g6486,g7906);
  and AND2_189(g8755,g3494,g8004);
  and AND2_190(g8760,g7053,g7845);
  and AND2_191(g8761,g7195,g8156);
  and AND2_192(g8762,g3806,g7892);
  and AND2_193(g8774,g6751,g7958);
  and AND2_194(g8778,g3650,g8079);
  and AND2_195(g8783,g7303,g7865);
  and AND2_196(g8784,g7391,g8242);
  and AND2_197(g8797,g7053,g8009);
  and AND2_198(g8801,g3806,g8164);
  and AND2_199(g8816,g7303,g8084);
  and AND2_200(g8841,g6486,g490);
  and AND2_201(g8842,g6512,g5508);
  and AND2_202(g8861,g6643,g493);
  and AND2_203(g8868,g6751,g1177);
  and AND2_204(g8869,g6776,g5552);
  and AND2_205(g8892,g3338,g496);
  and AND2_206(g8899,g6945,g1180);
  and AND2_207(g8906,g7053,g1871);
  and AND2_208(g8907,g7078,g5598);
  and AND2_209(g8932,g3494,g1183);
  and AND2_210(g8939,g7195,g1874);
  and AND2_211(g8946,g7303,g2565);
  and AND2_212(g8947,g7328,g5615);
  and AND2_213(g8972,g3650,g1877);
  and AND2_214(g8979,g7391,g2568);
  and AND2_215(g9004,g3806,g2571);
  and AND2_216(g9009,g6486,g565);
  and AND2_217(g9026,g5438,g7610);
  and AND2_218(g9033,g6643,g567);
  and AND2_219(g9034,g6751,g1251);
  and AND2_220(g9047,g6448,g7616);
  and AND2_221(g9048,g3338,g489);
  and AND2_222(g9049,g5473,g7619);
  and AND2_223(g9056,g6945,g1253);
  and AND2_224(g9057,g7053,g1945);
  and AND2_225(g9061,g3306,g7623);
  and AND2_226(g9062,g5438,g7626);
  and AND2_227(g9063,g5438,g7629);
  and AND2_228(g9064,g6713,g7632);
  and AND2_229(g9065,g3494,g1176);
  and AND2_230(g9066,g5512,g7635);
  and AND2_231(g9073,g7195,g1947);
  and AND2_232(g9074,g7303,g2639);
  and AND2_233(g9075,g6448,g7643);
  and AND2_234(g9076,g5438,g7646);
  and AND2_235(g9077,g6448,g7649);
  and AND2_236(g9078,g3462,g7652);
  and AND2_237(g9079,g5473,g7655);
  and AND2_238(g9080,g5473,g7658);
  and AND2_239(g9081,g7015,g7661);
  and AND2_240(g9082,g3650,g1870);
  and AND2_241(g9083,g5556,g7664);
  and AND2_242(g9090,g7391,g2641);
  and AND2_243(g9091,g3306,g7670);
  and AND2_244(g9092,g6448,g7673);
  and AND2_245(g9093,g3306,g7676);
  and AND2_246(g9094,g6713,g7679);
  and AND2_247(g9095,g5473,g7682);
  and AND2_248(g9096,g6713,g7685);
  and AND2_249(g9097,g3618,g7688);
  and AND2_250(g9098,g5512,g7691);
  and AND2_251(g9099,g5512,g7694);
  and AND2_252(g9100,g7265,g7697);
  and AND2_253(g9101,g3806,g2564);
  and AND2_254(g9102,g3306,g7703);
  and AND2_255(g9103,g3462,g7706);
  and AND2_256(g9104,g6713,g7709);
  and AND2_257(g9105,g3462,g7712);
  and AND2_258(g9106,g7015,g7715);
  and AND2_259(g9107,g5512,g7718);
  and AND2_260(g9108,g7015,g7721);
  and AND2_261(g9109,g3774,g7724);
  and AND2_262(g9110,g5556,g7727);
  and AND2_263(g9111,g5556,g7730);
  and AND2_264(g9112,g3462,g7733);
  and AND2_265(g9113,g3618,g7736);
  and AND2_266(g9114,g7015,g7739);
  and AND2_267(g9115,g3618,g7742);
  and AND2_268(g9116,g7265,g7745);
  and AND2_269(g9117,g5556,g7748);
  and AND2_270(g9118,g7265,g7751);
  and AND2_271(g9119,g5438,g7754);
  and AND2_272(g9120,g3618,g7757);
  and AND2_273(g9121,g3774,g7760);
  and AND2_274(g9122,g7265,g7763);
  and AND2_275(g9123,g3774,g7766);
  and AND2_276(g9124,g6448,g7769);
  and AND2_277(g9125,g5473,g7776);
  and AND2_278(g9126,g3774,g7779);
  and AND2_279(g9127,g3306,g7782);
  and AND2_280(g9131,g6713,g7785);
  and AND2_281(g9132,g5512,g7792);
  and AND2_282(g9133,g3462,g7796);
  and AND2_283(g9137,g7015,g7799);
  and AND2_284(g9138,g5556,g7806);
  and AND2_285(g9139,g3618,g7809);
  and AND2_286(g9143,g7265,g7812);
  and AND2_287(g9145,g3774,g7823);
  and AND2_288(g9241,g6232,g7950);
  and AND2_289(g9301,g6314,g7990);
  and AND2_290(g9302,g6232,g7993);
  and AND2_291(g9319,g6369,g8001);
  and AND2_292(g9364,g3254,g8053);
  and AND2_293(g9365,g6314,g8056);
  and AND2_294(g9366,g6232,g8059);
  and AND2_295(g9367,g6232,g8062);
  and AND2_296(g9382,g6519,g8065);
  and AND2_297(g9383,g6369,g8068);
  and AND2_298(g9400,g6574,g8076);
  and AND2_299(g9438,g3254,g8123);
  and AND2_300(g9439,g6314,g8126);
  and AND2_301(g9440,g6232,g8129);
  and AND2_302(g9441,g6314,g8132);
  and AND2_303(g9442,g6232,g8135);
  and AND2_304(g9461,g3410,g8138);
  and AND2_305(g9462,g6519,g8141);
  and AND2_306(g9463,g6369,g8144);
  and AND2_307(g9464,g6369,g8147);
  and AND2_308(g9479,g6783,g8150);
  and AND2_309(g9480,g6574,g8153);
  and AND2_310(g9497,g6838,g8161);
  and AND2_311(g9518,g3254,g8191);
  and AND2_312(g9519,g6314,g8194);
  and AND2_313(g9520,g6232,g8197);
  and AND2_314(g9521,g3254,g8200);
  and AND2_315(g9522,g6314,g8203);
  and AND2_316(g9523,g6232,g8206);
  and AND3_0(g9534,g7772,g6135,g538);
  and AND2_317(g9580,g3410,g8209);
  and AND2_318(g9581,g6519,g8212);
  and AND2_319(g9582,g6369,g8215);
  and AND2_320(g9583,g6519,g8218);
  and AND2_321(g9584,g6369,g8221);
  and AND2_322(g9603,g3566,g8224);
  and AND2_323(g9604,g6783,g8227);
  and AND2_324(g9605,g6574,g8230);
  and AND2_325(g9606,g6574,g8233);
  and AND2_326(g9621,g7085,g8236);
  and AND2_327(g9622,g6838,g8239);
  and AND2_328(g9630,g3254,g3922);
  and AND2_329(g9631,g6314,g3925);
  and AND2_330(g9632,g6232,g3928);
  and AND2_331(g9633,g3254,g3931);
  and AND2_332(g9634,g6314,g3934);
  and AND2_333(g9635,g6232,g3937);
  and AND4_0(II16735,g5856,g4338,g4339,g5141);
  and AND4_1(II16736,g5713,g5958,g4735,g4736);
  and AND2_334(g9636,II16735,II16736);
  and AND2_335(g9639,g5438,g408);
  and AND2_336(g9647,g6678,g3942);
  and AND2_337(g9648,g6678,g3945);
  and AND2_338(g9660,g3410,g3948);
  and AND2_339(g9661,g6519,g3951);
  and AND2_340(g9662,g6369,g3954);
  and AND2_341(g9663,g3410,g3957);
  and AND2_342(g9664,g6519,g3960);
  and AND2_343(g9665,g6369,g3963);
  and AND3_1(g9676,g7788,g6145,g1224);
  and AND2_344(g9722,g3566,g3966);
  and AND2_345(g9723,g6783,g3969);
  and AND2_346(g9724,g6574,g3972);
  and AND2_347(g9725,g6783,g3975);
  and AND2_348(g9726,g6574,g3978);
  and AND2_349(g9745,g3722,g3981);
  and AND2_350(g9746,g7085,g3984);
  and AND2_351(g9747,g6838,g3987);
  and AND2_352(g9748,g6838,g3990);
  and AND2_353(g9759,g3254,g4000);
  and AND2_354(g9760,g6314,g4003);
  and AND2_355(g9761,g6232,g4006);
  and AND2_356(g9762,g3254,g4009);
  and AND2_357(g9763,g6314,g4012);
  and AND2_358(g9764,g6448,g411);
  and AND2_359(g9765,g5438,g417);
  and AND2_360(g9766,g5438,g4017);
  and AND2_361(g9773,g6912,g4020);
  and AND2_362(g9774,g6678,g4023);
  and AND2_363(g9775,g6912,g4026);
  and AND2_364(g9776,g3410,g4029);
  and AND2_365(g9777,g6519,g4032);
  and AND2_366(g9778,g6369,g4035);
  and AND2_367(g9779,g3410,g4038);
  and AND2_368(g9780,g6519,g4041);
  and AND2_369(g9781,g6369,g4044);
  and AND4_2(II16826,g5903,g4507,g4508,g5234);
  and AND4_3(II16827,g5771,g5987,g4911,g4912);
  and AND2_370(g9782,II16826,II16827);
  and AND2_371(g9785,g5473,g1095);
  and AND2_372(g9793,g6980,g4049);
  and AND2_373(g9794,g6980,g4052);
  and AND2_374(g9806,g3566,g4055);
  and AND2_375(g9807,g6783,g4058);
  and AND2_376(g9808,g6574,g4061);
  and AND2_377(g9809,g3566,g4064);
  and AND2_378(g9810,g6783,g4067);
  and AND2_379(g9811,g6574,g4070);
  and AND3_2(g9822,g7802,g6166,g1918);
  and AND2_380(g9868,g3722,g4073);
  and AND2_381(g9869,g7085,g4076);
  and AND2_382(g9870,g6838,g4079);
  and AND2_383(g9871,g7085,g4082);
  and AND2_384(g9872,g6838,g4085);
  and AND2_385(g9887,g6232,g4095);
  and AND2_386(g9888,g3254,g4098);
  and AND2_387(g9889,g6314,g4101);
  and AND2_388(g9890,g6232,g4104);
  and AND2_389(g9891,g3254,g4107);
  and AND2_390(g9892,g3306,g414);
  and AND2_391(g9893,g6448,g420);
  and AND2_392(g9894,g6448,g4112);
  and AND2_393(g9901,g3366,g4115);
  and AND2_394(g9902,g6912,g4118);
  and AND2_395(g9903,g6678,g4121);
  and AND2_396(g9904,g3366,g4124);
  and AND2_397(g9905,g3410,g4127);
  and AND2_398(g9906,g6519,g4130);
  and AND2_399(g9907,g6369,g4133);
  and AND2_400(g9908,g3410,g4136);
  and AND2_401(g9909,g6519,g4139);
  and AND2_402(g9910,g6713,g1098);
  and AND2_403(g9911,g5473,g1104);
  and AND2_404(g9912,g5473,g4144);
  and AND2_405(g9919,g7162,g4147);
  and AND2_406(g9920,g6980,g4150);
  and AND2_407(g9921,g7162,g4153);
  and AND2_408(g9922,g3566,g4156);
  and AND2_409(g9923,g6783,g4159);
  and AND2_410(g9924,g6574,g4162);
  and AND2_411(g9925,g3566,g4165);
  and AND2_412(g9926,g6783,g4168);
  and AND2_413(g9927,g6574,g4171);
  and AND4_4(II16930,g5942,g4683,g4684,g5297);
  and AND4_5(II16931,g5830,g6024,g5070,g5071);
  and AND2_414(g9928,II16930,II16931);
  and AND2_415(g9931,g5512,g1789);
  and AND2_416(g9939,g7230,g4176);
  and AND2_417(g9940,g7230,g4179);
  and AND2_418(g9952,g3722,g4182);
  and AND2_419(g9953,g7085,g4185);
  and AND2_420(g9954,g6838,g4188);
  and AND2_421(g9955,g3722,g4191);
  and AND2_422(g9956,g7085,g4194);
  and AND2_423(g9957,g6838,g4197);
  and AND3_3(g9968,g7815,g6193,g2612);
  and AND2_424(g10007,g6314,g4205);
  and AND2_425(g10008,g6232,g4208);
  and AND2_426(g10009,g3254,g4211);
  and AND2_427(g10010,g6314,g4214);
  and AND2_428(g10011,g5438,g4217);
  and AND2_429(g10012,g3306,g423);
  and AND2_430(g10013,g3306,g4221);
  and AND2_431(g10014,g5438,g429);
  and AND2_432(g10024,g3398,g6912);
  and AND2_433(g10035,g3366,g4225);
  and AND2_434(g10036,g6912,g4228);
  and AND2_435(g10037,g6678,g4231);
  and AND2_436(g10041,g6369,g4234);
  and AND2_437(g10042,g3410,g4237);
  and AND2_438(g10043,g6519,g4240);
  and AND2_439(g10044,g6369,g4243);
  and AND2_440(g10045,g3410,g4246);
  and AND2_441(g10046,g3462,g1101);
  and AND2_442(g10047,g6713,g1107);
  and AND2_443(g10048,g6713,g4251);
  and AND2_444(g10055,g3522,g4254);
  and AND2_445(g10056,g7162,g4257);
  and AND2_446(g10057,g6980,g4260);
  and AND2_447(g10058,g3522,g4263);
  and AND2_448(g10059,g3566,g4266);
  and AND2_449(g10060,g6783,g4269);
  and AND2_450(g10061,g6574,g4272);
  and AND2_451(g10062,g3566,g4275);
  and AND2_452(g10063,g6783,g4278);
  and AND2_453(g10064,g7015,g1792);
  and AND2_454(g10065,g5512,g1798);
  and AND2_455(g10066,g5512,g4283);
  and AND2_456(g10073,g7358,g4286);
  and AND2_457(g10074,g7230,g4289);
  and AND2_458(g10075,g7358,g4292);
  and AND2_459(g10076,g3722,g4295);
  and AND2_460(g10077,g7085,g4298);
  and AND2_461(g10078,g6838,g4301);
  and AND2_462(g10079,g3722,g4304);
  and AND2_463(g10080,g7085,g4307);
  and AND2_464(g10081,g6838,g4310);
  and AND4_6(II17042,g5976,g4860,g4861,g5334);
  and AND4_7(II17043,g5886,g6040,g5199,g5200);
  and AND2_465(g10082,II17042,II17043);
  and AND2_466(g10085,g5556,g2483);
  and AND2_467(g10093,g7426,g4315);
  and AND2_468(g10094,g7426,g4318);
  and AND2_469(g10101,g3254,g4329);
  and AND2_470(g10102,g6314,g4332);
  and AND2_471(g10103,g3254,g4335);
  and AND2_472(g10104,g6448,g4340);
  and AND2_473(g10105,g5438,g4343);
  and AND2_474(g10106,g6448,g432);
  and AND2_475(g10107,g5438,g438);
  and AND2_476(g10108,g6486,g569);
  and AND2_477(g10112,g3366,g4348);
  and AND2_478(g10113,g6912,g4351);
  and AND2_479(g10114,g6678,g4354);
  and AND2_480(g10115,g6678,g4357);
  and AND2_481(g10116,g6519,g4360);
  and AND2_482(g10117,g6369,g4363);
  and AND2_483(g10118,g3410,g4366);
  and AND2_484(g10119,g6519,g4369);
  and AND2_485(g10120,g5473,g4372);
  and AND2_486(g10121,g3462,g1110);
  and AND2_487(g10122,g3462,g4376);
  and AND2_488(g10123,g5473,g1116);
  and AND2_489(g10133,g3554,g7162);
  and AND2_490(g10144,g3522,g4380);
  and AND2_491(g10145,g7162,g4383);
  and AND2_492(g10146,g6980,g4386);
  and AND2_493(g10150,g6574,g4389);
  and AND2_494(g10151,g3566,g4392);
  and AND2_495(g10152,g6783,g4395);
  and AND2_496(g10153,g6574,g4398);
  and AND2_497(g10154,g3566,g4401);
  and AND2_498(g10155,g3618,g1795);
  and AND2_499(g10156,g7015,g1801);
  and AND2_500(g10157,g7015,g4406);
  and AND2_501(g10164,g3678,g4409);
  and AND2_502(g10165,g7358,g4412);
  and AND2_503(g10166,g7230,g4415);
  and AND2_504(g10167,g3678,g4418);
  and AND2_505(g10168,g3722,g4421);
  and AND2_506(g10169,g7085,g4424);
  and AND2_507(g10170,g6838,g4427);
  and AND2_508(g10171,g3722,g4430);
  and AND2_509(g10172,g7085,g4433);
  and AND2_510(g10173,g7265,g2486);
  and AND2_511(g10174,g5556,g2492);
  and AND2_512(g10175,g5556,g4438);
  and AND2_513(g10182,g7488,g4441);
  and AND2_514(g10183,g7426,g4444);
  and AND2_515(g10184,g7488,g4447);
  and AND4_8(II17156,g6898,g2998,g6901,g3002);
  and AND4_9(g10186,g3013,g7466,g3024,II17156);
  and AND2_516(g10192,g3254,g4453);
  and AND2_517(g10193,g3306,g4465);
  and AND2_518(g10194,g6448,g4468);
  and AND2_519(g10195,g5438,g4471);
  and AND2_520(g10196,g3306,g435);
  and AND2_521(g10197,g6448,g441);
  and AND2_522(g10198,g6643,g571);
  and AND2_523(g10199,g6486,g4476);
  and AND2_524(g10200,g6486,g587);
  and AND2_525(g10201,g3366,g4480);
  and AND2_526(g10202,g6912,g4483);
  and AND2_527(g10203,g6678,g4486);
  and AND2_528(g10204,g6912,g4489);
  and AND2_529(g10205,g6678,g4492);
  and AND2_530(g10206,g3410,g4498);
  and AND2_531(g10207,g6519,g4501);
  and AND2_532(g10208,g3410,g4504);
  and AND2_533(g10209,g6713,g4509);
  and AND2_534(g10210,g5473,g4512);
  and AND2_535(g10211,g6713,g1119);
  and AND2_536(g10212,g5473,g1125);
  and AND2_537(g10213,g6751,g1255);
  and AND2_538(g10217,g3522,g4517);
  and AND2_539(g10218,g7162,g4520);
  and AND2_540(g10219,g6980,g4523);
  and AND2_541(g10220,g6980,g4526);
  and AND2_542(g10221,g6783,g4529);
  and AND2_543(g10222,g6574,g4532);
  and AND2_544(g10223,g3566,g4535);
  and AND2_545(g10224,g6783,g4538);
  and AND2_546(g10225,g5512,g4541);
  and AND2_547(g10226,g3618,g1804);
  and AND2_548(g10227,g3618,g4545);
  and AND2_549(g10228,g5512,g1810);
  and AND2_550(g10238,g3710,g7358);
  and AND2_551(g10249,g3678,g4549);
  and AND2_552(g10250,g7358,g4552);
  and AND2_553(g10251,g7230,g4555);
  and AND2_554(g10255,g6838,g4558);
  and AND2_555(g10256,g3722,g4561);
  and AND2_556(g10257,g7085,g4564);
  and AND2_557(g10258,g6838,g4567);
  and AND2_558(g10259,g3722,g4570);
  and AND2_559(g10260,g3774,g2489);
  and AND2_560(g10261,g7265,g2495);
  and AND2_561(g10262,g7265,g4575);
  and AND2_562(g10269,g3834,g4578);
  and AND2_563(g10270,g7488,g4581);
  and AND2_564(g10271,g7426,g4584);
  and AND2_565(g10272,g3834,g4587);
  and AND2_566(g10279,g3306,g4592);
  and AND2_567(g10280,g6448,g4595);
  and AND2_568(g10281,g5438,g4598);
  and AND2_569(g10282,g3306,g444);
  and AND2_570(g10283,g3338,g573);
  and AND2_571(g10284,g6643,g4603);
  and AND2_572(g10285,g6486,g4606);
  and AND2_573(g10286,g6643,g590);
  and AND2_574(g10287,g6486,g596);
  and AND2_575(g10288,g3366,g4611);
  and AND2_576(g10289,g6912,g4614);
  and AND2_577(g10290,g6678,g4617);
  and AND2_578(g10291,g3366,g4620);
  and AND2_579(g10292,g6912,g4623);
  and AND2_580(g10293,g6678,g4626);
  and AND2_581(g10294,g3410,g4629);
  and AND2_582(g10295,g3462,g4641);
  and AND2_583(g10296,g6713,g4644);
  and AND2_584(g10297,g5473,g4647);
  and AND2_585(g10298,g3462,g1122);
  and AND2_586(g10299,g6713,g1128);
  and AND2_587(g10300,g6945,g1257);
  and AND2_588(g10301,g6751,g4652);
  and AND2_589(g10302,g6751,g1273);
  and AND2_590(g10303,g3522,g4656);
  and AND2_591(g10304,g7162,g4659);
  and AND2_592(g10305,g6980,g4662);
  and AND2_593(g10306,g7162,g4665);
  and AND2_594(g10307,g6980,g4668);
  and AND2_595(g10308,g3566,g4674);
  and AND2_596(g10309,g6783,g4677);
  and AND2_597(g10310,g3566,g4680);
  and AND2_598(g10311,g7015,g4685);
  and AND2_599(g10312,g5512,g4688);
  and AND2_600(g10313,g7015,g1813);
  and AND2_601(g10314,g5512,g1819);
  and AND2_602(g10315,g7053,g1949);
  and AND2_603(g10319,g3678,g4693);
  and AND2_604(g10320,g7358,g4696);
  and AND2_605(g10321,g7230,g4699);
  and AND2_606(g10322,g7230,g4702);
  and AND2_607(g10323,g7085,g4705);
  and AND2_608(g10324,g6838,g4708);
  and AND2_609(g10325,g3722,g4711);
  and AND2_610(g10326,g7085,g4714);
  and AND2_611(g10327,g5556,g4717);
  and AND2_612(g10328,g3774,g2498);
  and AND2_613(g10329,g3774,g4721);
  and AND2_614(g10330,g5556,g2504);
  and AND2_615(g10340,g3866,g7488);
  and AND2_616(g10351,g3834,g4725);
  and AND2_617(g10352,g7488,g4728);
  and AND2_618(g10353,g7426,g4731);
  and AND2_619(g10360,g3306,g4737);
  and AND2_620(g10361,g6448,g4740);
  and AND2_621(g10362,g3338,g4743);
  and AND2_622(g10363,g6643,g4746);
  and AND2_623(g10364,g6486,g4749);
  and AND2_624(g10365,g3338,g593);
  and AND2_625(g10366,g6643,g599);
  and AND2_626(g10367,g3366,g4754);
  and AND2_627(g10368,g6912,g4757);
  and AND2_628(g10369,g6678,g4760);
  and AND2_629(g10370,g3366,g4763);
  and AND2_630(g10371,g6912,g4766);
  and AND2_631(g10372,g3462,g4769);
  and AND2_632(g10373,g6713,g4772);
  and AND2_633(g10374,g5473,g4775);
  and AND2_634(g10375,g3462,g1131);
  and AND2_635(g10376,g3494,g1259);
  and AND2_636(g10377,g6945,g4780);
  and AND2_637(g10378,g6751,g4783);
  and AND2_638(g10379,g6945,g1276);
  and AND2_639(g10380,g6751,g1282);
  and AND2_640(g10381,g3522,g4788);
  and AND2_641(g10382,g7162,g4791);
  and AND2_642(g10383,g6980,g4794);
  and AND2_643(g10384,g3522,g4797);
  and AND2_644(g10385,g7162,g4800);
  and AND2_645(g10386,g6980,g4803);
  and AND2_646(g10387,g3566,g4806);
  and AND2_647(g10388,g3618,g4818);
  and AND2_648(g10389,g7015,g4821);
  and AND2_649(g10390,g5512,g4824);
  and AND2_650(g10391,g3618,g1816);
  and AND2_651(g10392,g7015,g1822);
  and AND2_652(g10393,g7195,g1951);
  and AND2_653(g10394,g7053,g4829);
  and AND2_654(g10395,g7053,g1967);
  and AND2_655(g10396,g3678,g4833);
  and AND2_656(g10397,g7358,g4836);
  and AND2_657(g10398,g7230,g4839);
  and AND2_658(g10399,g7358,g4842);
  and AND2_659(g10400,g7230,g4845);
  and AND2_660(g10401,g3722,g4851);
  and AND2_661(g10402,g7085,g4854);
  and AND2_662(g10403,g3722,g4857);
  and AND2_663(g10404,g7265,g4862);
  and AND2_664(g10405,g5556,g4865);
  and AND2_665(g10406,g7265,g2507);
  and AND2_666(g10407,g5556,g2513);
  and AND2_667(g10408,g7303,g2643);
  and AND2_668(g10412,g3834,g4870);
  and AND2_669(g10413,g7488,g4873);
  and AND2_670(g10414,g7426,g4876);
  and AND2_671(g10415,g7426,g4879);
  and AND2_672(g10422,g3306,g4882);
  and AND2_673(g10423,g5438,g4885);
  and AND2_674(g10430,g3338,g4888);
  and AND2_675(g10431,g6643,g4891);
  and AND2_676(g10432,g6486,g4894);
  and AND2_677(g10433,g3338,g602);
  and AND2_678(g10434,g6486,g605);
  and AND2_679(g10435,g3366,g4899);
  and AND2_680(g10436,g6912,g4902);
  and AND2_681(g10437,g6678,g4905);
  and AND2_682(g10438,g3366,g4908);
  and AND2_683(g10439,g3462,g4913);
  and AND2_684(g10440,g6713,g4916);
  and AND2_685(g10441,g3494,g4919);
  and AND2_686(g10442,g6945,g4922);
  and AND2_687(g10443,g6751,g4925);
  and AND2_688(g10444,g3494,g1279);
  and AND2_689(g10445,g6945,g1285);
  and AND2_690(g10446,g3522,g4930);
  and AND2_691(g10447,g7162,g4933);
  and AND2_692(g10448,g6980,g4936);
  and AND2_693(g10449,g3522,g4939);
  and AND2_694(g10450,g7162,g4942);
  and AND2_695(g10451,g3618,g4945);
  and AND2_696(g10452,g7015,g4948);
  and AND2_697(g10453,g5512,g4951);
  and AND2_698(g10454,g3618,g1825);
  and AND2_699(g10455,g3650,g1953);
  and AND2_700(g10456,g7195,g4956);
  and AND2_701(g10457,g7053,g4959);
  and AND2_702(g10458,g7195,g1970);
  and AND2_703(g10459,g7053,g1976);
  and AND2_704(g10460,g3678,g4964);
  and AND2_705(g10461,g7358,g4967);
  and AND2_706(g10462,g7230,g4970);
  and AND2_707(g10463,g3678,g4973);
  and AND2_708(g10464,g7358,g4976);
  and AND2_709(g10465,g7230,g4979);
  and AND2_710(g10466,g3722,g4982);
  and AND2_711(g10467,g3774,g4994);
  and AND2_712(g10468,g7265,g4997);
  and AND2_713(g10469,g5556,g5000);
  and AND2_714(g10470,g3774,g2510);
  and AND2_715(g10471,g7265,g2516);
  and AND2_716(g10472,g7391,g2645);
  and AND2_717(g10473,g7303,g5005);
  and AND2_718(g10474,g7303,g2661);
  and AND2_719(g10475,g3834,g5009);
  and AND2_720(g10476,g7488,g5012);
  and AND2_721(g10477,g7426,g5015);
  and AND2_722(g10478,g7488,g5018);
  and AND2_723(g10479,g7426,g5021);
  and AND3_4(II17429,g6901,g7338,g7146);
  and AND3_5(g10480,g7466,g7342,II17429);
  and AND2_724(g10485,g6448,g5024);
  and AND2_725(g10492,g3338,g5027);
  and AND2_726(g10493,g6643,g5030);
  and AND2_727(g10494,g6643,g608);
  and AND2_728(g10495,g6486,g614);
  and AND2_729(g10496,g3366,g5035);
  and AND2_730(g10497,g6912,g5038);
  and AND2_731(g10498,g3462,g5041);
  and AND2_732(g10499,g5473,g5044);
  and AND2_733(g10506,g3494,g5047);
  and AND2_734(g10507,g6945,g5050);
  and AND2_735(g10508,g6751,g5053);
  and AND2_736(g10509,g3494,g1288);
  and AND2_737(g10510,g6751,g1291);
  and AND2_738(g10511,g3522,g5058);
  and AND2_739(g10512,g7162,g5061);
  and AND2_740(g10513,g6980,g5064);
  and AND2_741(g10514,g3522,g5067);
  and AND2_742(g10515,g3618,g5072);
  and AND2_743(g10516,g7015,g5075);
  and AND2_744(g10517,g3650,g5078);
  and AND2_745(g10518,g7195,g5081);
  and AND2_746(g10519,g7053,g5084);
  and AND2_747(g10520,g3650,g1973);
  and AND2_748(g10521,g7195,g1979);
  and AND2_749(g10522,g3678,g5089);
  and AND2_750(g10523,g7358,g5092);
  and AND2_751(g10524,g7230,g5095);
  and AND2_752(g10525,g3678,g5098);
  and AND2_753(g10526,g7358,g5101);
  and AND2_754(g10527,g3774,g5104);
  and AND2_755(g10528,g7265,g5107);
  and AND2_756(g10529,g5556,g5110);
  and AND2_757(g10530,g3774,g2519);
  and AND2_758(g10531,g3806,g2647);
  and AND2_759(g10532,g7391,g5115);
  and AND2_760(g10533,g7303,g5118);
  and AND2_761(g10534,g7391,g2664);
  and AND2_762(g10535,g7303,g2670);
  and AND2_763(g10536,g3834,g5123);
  and AND2_764(g10537,g7488,g5126);
  and AND2_765(g10538,g7426,g5129);
  and AND2_766(g10539,g3834,g5132);
  and AND2_767(g10540,g7488,g5135);
  and AND2_768(g10541,g7426,g5138);
  and AND2_769(g10548,g3306,g5142);
  and AND2_770(g10555,g3338,g5145);
  and AND2_771(g10556,g3338,g611);
  and AND2_772(g10557,g6643,g617);
  and AND2_773(g10558,g3366,g5150);
  and AND2_774(g10559,g6713,g5153);
  and AND2_775(g10566,g3494,g5156);
  and AND2_776(g10567,g6945,g5159);
  and AND2_777(g10568,g6945,g1294);
  and AND2_778(g10569,g6751,g1300);
  and AND2_779(g10570,g3522,g5164);
  and AND2_780(g10571,g7162,g5167);
  and AND2_781(g10572,g3618,g5170);
  and AND2_782(g10573,g5512,g5173);
  and AND2_783(g10580,g3650,g5176);
  and AND2_784(g10581,g7195,g5179);
  and AND2_785(g10582,g7053,g5182);
  and AND2_786(g10583,g3650,g1982);
  and AND2_787(g10584,g7053,g1985);
  and AND2_788(g10585,g3678,g5187);
  and AND2_789(g10586,g7358,g5190);
  and AND2_790(g10587,g7230,g5193);
  and AND2_791(g10588,g3678,g5196);
  and AND2_792(g10589,g3774,g5201);
  and AND2_793(g10590,g7265,g5204);
  and AND2_794(g10591,g3806,g5207);
  and AND2_795(g10592,g7391,g5210);
  and AND2_796(g10593,g7303,g5213);
  and AND2_797(g10594,g3806,g2667);
  and AND2_798(g10595,g7391,g2673);
  and AND2_799(g10596,g3834,g5218);
  and AND2_800(g10597,g7488,g5221);
  and AND2_801(g10598,g7426,g5224);
  and AND2_802(g10599,g3834,g5227);
  and AND2_803(g10600,g7488,g5230);
  and AND2_804(g10604,g3338,g620);
  and AND2_805(g10605,g3462,g5235);
  and AND2_806(g10612,g3494,g5238);
  and AND2_807(g10613,g3494,g1297);
  and AND2_808(g10614,g6945,g1303);
  and AND2_809(g10615,g3522,g5243);
  and AND2_810(g10616,g7015,g5246);
  and AND2_811(g10623,g3650,g5249);
  and AND2_812(g10624,g7195,g5252);
  and AND2_813(g10625,g7195,g1988);
  and AND2_814(g10626,g7053,g1994);
  and AND2_815(g10627,g3678,g5257);
  and AND2_816(g10628,g7358,g5260);
  and AND2_817(g10629,g3774,g5263);
  and AND2_818(g10630,g5556,g5266);
  and AND2_819(g10637,g3806,g5269);
  and AND2_820(g10638,g7391,g5272);
  and AND2_821(g10639,g7303,g5275);
  and AND2_822(g10640,g3806,g2676);
  and AND2_823(g10641,g7303,g2679);
  and AND2_824(g10642,g3834,g5280);
  and AND2_825(g10643,g7488,g5283);
  and AND2_826(g10644,g7426,g5286);
  and AND2_827(g10645,g3834,g5289);
  and AND2_828(g10650,g6678,g5293);
  and AND2_829(g10651,g3494,g1306);
  and AND2_830(g10652,g3618,g5298);
  and AND2_831(g10659,g3650,g5301);
  and AND2_832(g10660,g3650,g1991);
  and AND2_833(g10661,g7195,g1997);
  and AND2_834(g10662,g3678,g5306);
  and AND2_835(g10663,g7265,g5309);
  and AND2_836(g10670,g3806,g5312);
  and AND2_837(g10671,g7391,g5315);
  and AND2_838(g10672,g7391,g2682);
  and AND2_839(g10673,g7303,g2688);
  and AND2_840(g10674,g3834,g5320);
  and AND2_841(g10675,g7488,g5323);
  and AND2_842(g10678,g6912,g5327);
  and AND2_843(g10680,g6980,g5330);
  and AND2_844(g10681,g3650,g2000);
  and AND2_845(g10682,g3774,g5335);
  and AND2_846(g10689,g3806,g5338);
  and AND2_847(g10690,g3806,g2685);
  and AND2_848(g10691,g7391,g2691);
  and AND2_849(g10692,g3834,g5343);
  and AND4_10(g10693,g7462,g7522,g2924,g7545);
  and AND2_850(g10704,g3366,g5352);
  and AND2_851(g10707,g7162,g5355);
  and AND2_852(g10709,g7230,g5358);
  and AND2_853(g10710,g3806,g2694);
  and AND3_6(II17599,g7566,g7583,g7587);
  and AND3_7(g10711,g7595,g7600,II17599);
  and AND2_854(g10724,g3522,g5369);
  and AND2_855(g10727,g7358,g5372);
  and AND2_856(g10729,g7426,g5375);
  and AND2_857(g10745,g3678,g5382);
  and AND2_858(g10748,g7488,g5385);
  and AND2_859(g10764,g3834,g5391);
  and AND2_860(g11347,g6232,g213);
  and AND2_861(g11420,g6314,g216);
  and AND2_862(g11421,g6232,g222);
  and AND2_863(g11431,g6369,g900);
  and AND2_864(g11607,g5871,g8360);
  and AND2_865(g11612,g5881,g8378);
  and AND2_866(g11637,g5918,g8427);
  and AND2_867(g11771,g554,g8622);
  and AND2_868(g11788,g1240,g8632);
  and AND2_869(g11805,g6173,g8643);
  and AND2_870(g11814,g1934,g8651);
  and AND2_871(g11816,g7869,g8655);
  and AND2_872(g11838,g6205,g8659);
  and AND2_873(g11847,g2628,g8667);
  and AND2_874(g11851,g7849,g8670);
  and AND2_875(g11880,g6294,g8678);
  and AND2_876(g11885,g7834,g8684);
  and AND2_877(g11922,g6431,g8690);
  and AND2_878(g11926,g8169,g8696);
  and AND2_879(g11966,g8090,g8708);
  and AND2_880(g11967,g7967,g8711);
  and AND2_881(g12012,g8015,g8745);
  and AND2_882(g12069,g7964,g8763);
  and AND2_883(g12070,g8018,g8766);
  and AND2_884(g12128,g7916,g8785);
  and AND2_885(g12129,g7872,g8788);
  and AND2_886(g12186,g8093,g8805);
  and AND2_887(g12273,g8172,g8829);
  and AND2_888(g12274,g7900,g8832);
  and AND2_889(g12307,g7919,g8853);
  and AND2_890(g12330,g8246,g8879);
  and AND2_891(g12331,g7927,g8882);
  and AND2_892(g12353,g7852,g8915);
  and AND2_893(g12376,g7974,g8949);
  and AND2_894(g12419,g8028,g9006);
  and AND2_895(g12429,g8101,g9044);
  and AND2_896(g12477,g7822,g9128);
  and AND2_897(g12494,g7833,g9134);
  and AND2_898(g12514,g7848,g9140);
  and AND2_899(g12531,g7868,g9146);
  and AND2_900(g12650,g6149,g9290);
  and AND4_11(II19937,g9507,g9427,g9356,g9293);
  and AND4_12(II19938,g9232,g9187,g9161,g9150);
  and AND2_901(g12876,II19937,II19938);
  and AND2_902(g12908,g7899,g10004);
  and AND4_13(II19971,g9649,g9569,g9453,g9374);
  and AND4_14(II19972,g9310,g9248,g9203,g9174);
  and AND2_903(g12916,II19971,II19972);
  and AND2_904(g12938,g8179,g10096);
  and AND4_15(II19996,g9795,g9711,g9595,g9471);
  and AND4_16(II19997,g9391,g9326,g9264,g9216);
  and AND2_905(g12945,II19996,II19997);
  and AND2_906(g12966,g7926,g10189);
  and AND4_17(II20021,g9941,g9857,g9737,g9613);
  and AND4_18(II20022,g9488,g9407,g9342,g9277);
  and AND2_907(g12974,II20021,II20022);
  and AND2_908(g12989,g8254,g10273);
  and AND2_909(g12990,g8180,g10276);
  and AND2_910(g13000,g7973,g10357);
  and AND2_911(g13004,g10186,g8317);
  and AND2_912(g13009,g3995,g10416);
  and AND2_913(g13010,g8255,g10419);
  and AND2_914(g13023,g8027,g10482);
  and AND2_915(g13031,g7879,g10542);
  and AND2_916(g13032,g3996,g10545);
  and AND2_917(g13042,g8100,g10601);
  and AND3_8(II20100,g10186,g3018,g3028);
  and AND3_9(g13055,g7471,g7570,II20100);
  and AND2_918(g13056,g4092,g10646);
  and AND4_19(II20131,g8313,g7542,g2888,g7566);
  and AND4_20(II20132,g2892,g2903,g7595,g2908);
  and AND2_919(g13082,II20131,II20132);
  and AND4_21(g13110,g10693,g2883,g7562,g10711);
  and AND2_920(g13247,g298,g11032);
  and AND2_921(g13266,g5628,g11088);
  and AND2_922(g13270,g985,g11102);
  and AND2_923(g13289,g5647,g11141);
  and AND2_924(g13291,g5656,g11154);
  and AND2_925(g13295,g1679,g11170);
  and AND2_926(g13316,g5675,g11210);
  and AND2_927(g13320,g5685,g11225);
  and AND2_928(g13322,g5694,g11240);
  and AND2_929(g13326,g2373,g11256);
  and AND2_930(g13335,g5708,g11278);
  and AND2_931(g13340,g5727,g11294);
  and AND2_932(g13343,g5737,g11309);
  and AND2_933(g13345,g5746,g11324);
  and AND2_934(g13355,g5756,g11355);
  and AND2_935(g13360,g5766,g11373);
  and AND2_936(g13365,g5785,g11389);
  and AND2_937(g13368,g5795,g11404);
  and AND2_938(g13385,g5815,g11441);
  and AND2_939(g13390,g5825,g11459);
  and AND2_940(g13395,g5844,g11475);
  and AND2_941(g13477,g6016,g12191);
  and AND2_942(g13479,g6017,g12196);
  and AND2_943(g13480,g6018,g12197);
  and AND2_944(g13481,g5864,g11603);
  and AND2_945(g13483,g6020,g12209);
  and AND2_946(g13484,g6021,g12210);
  and AND2_947(g13485,g6022,g12211);
  and AND2_948(g13486,g6023,g12212);
  and AND2_949(g13487,g5874,g11608);
  and AND2_950(g13488,g6025,g12218);
  and AND2_951(g13489,g6026,g12219);
  and AND2_952(g13490,g6027,g12220);
  and AND2_953(g13491,g6028,g12221);
  and AND2_954(g13492,g2371,g12222);
  and AND2_955(g13493,g5887,g11613);
  and AND2_956(g13496,g6032,g12246);
  and AND2_957(g13498,g6033,g12251);
  and AND2_958(g13499,g6034,g12252);
  and AND2_959(g13500,g5911,g11633);
  and AND2_960(g13502,g6036,g12264);
  and AND2_961(g13503,g6037,g12265);
  and AND2_962(g13504,g6038,g12266);
  and AND2_963(g13505,g6039,g12267);
  and AND2_964(g13506,g5921,g11638);
  and AND2_965(g13513,g6043,g12289);
  and AND2_966(g13515,g6044,g12294);
  and AND2_967(g13516,g6045,g12295);
  and AND2_968(g13517,g5950,g11656);
  and AND2_969(g13527,g6047,g12325);
  and AND2_970(g13609,g6141,g12456);
  and AND2_971(g13619,g6162,g12466);
  and AND2_972(g13623,g5428,g12472);
  and AND2_973(g13625,g6173,g12476);
  and AND2_974(g13631,g6189,g12481);
  and AND2_975(g13634,g12776,g8617);
  and AND2_976(g13636,g6205,g12493);
  and AND2_977(g13642,g6221,g12498);
  and AND2_978(g13643,g5431,g12502);
  and AND2_979(g13645,g6281,g12504);
  and AND2_980(g13646,g7772,g12505);
  and AND2_981(g13648,g6294,g12513);
  and AND2_982(g13654,g8093,g11791);
  and AND2_983(g13655,g7540,g12518);
  and AND2_984(g13656,g12776,g8640);
  and AND2_985(g13671,g6418,g12521);
  and AND2_986(g13672,g7788,g12522);
  and AND2_987(g13674,g6431,g12530);
  and AND2_988(g13675,g7561,g12532);
  and AND2_989(g13676,g5434,g12533);
  and AND2_990(g13701,g6623,g12536);
  and AND2_991(g13702,g7802,g12537);
  and AND2_992(g13703,g8018,g11848);
  and AND2_993(g13704,g7581,g12542);
  and AND2_994(g13705,g12776,g8673);
  and AND2_995(g13738,g6887,g12545);
  and AND2_996(g13739,g7815,g12546);
  and AND2_997(g13740,g6636,g12547);
  and AND2_998(g13755,g7347,g12551);
  and AND2_999(g13787,g7967,g11923);
  and AND2_1000(g13788,g6897,g12553);
  and AND2_1001(g13789,g7140,g12554);
  and AND2_1002(g13790,g7475,g12558);
  and AND2_1003(g13796,g7477,g12559);
  and AND2_1004(g13815,g7139,g12560);
  and AND2_1005(g13816,g7530,g12596);
  and AND2_1006(g13818,g7531,g12597);
  and AND2_1007(g13824,g7533,g12598);
  and AND2_1008(g13833,g7919,g12009);
  and AND2_1009(g13834,g7336,g12599);
  and AND2_1010(g13835,g7461,g12600);
  and AND2_1011(g13837,g7556,g12642);
  and AND2_1012(g13839,g7557,g12643);
  and AND2_1013(g13845,g7559,g12644);
  and AND2_1014(g13846,g7460,g12645);
  and AND2_1015(g13847,g7521,g12646);
  and AND2_1016(g13851,g7579,g12688);
  and AND2_1017(g13853,g7580,g12689);
  and AND2_1018(g13854,g5349,g12690);
  and AND2_1019(g13855,g7541,g12691);
  and AND2_1020(g13860,g7593,g12742);
  and AND2_1021(g13862,g5366,g12743);
  and AND2_1022(g13865,g548,g12748);
  and AND2_1023(g13870,g7582,g12768);
  and AND2_1024(g13871,g7898,g12775);
  and AND2_1025(g13878,g7610,g12782);
  and AND2_1026(g13880,g1234,g12790);
  and AND2_1027(g13884,g7594,g12807);
  and AND2_1028(g13892,g7616,g12815);
  and AND2_1029(g13900,g7619,g12821);
  and AND2_1030(g13902,g1928,g12829);
  and AND2_1031(g13904,g7337,g12843);
  and AND2_1032(g13905,g7925,g12847);
  and AND2_1033(g13913,g7623,g12850);
  and AND2_1034(g13914,g7626,g12851);
  and AND2_1035(g13933,g7632,g12853);
  and AND2_1036(g13941,g7635,g12859);
  and AND2_1037(g13943,g2622,g12867);
  and AND2_1038(g13944,g7141,g12874);
  and AND2_1039(g13952,g7643,g12881);
  and AND2_1040(g13953,g7646,g12882);
  and AND2_1041(g13969,g7652,g12891);
  and AND2_1042(g13970,g7655,g12892);
  and AND2_1043(g13989,g7661,g12894);
  and AND2_1044(g13997,g7664,g12900);
  and AND2_1045(g13998,g7972,g12907);
  and AND2_1046(g14006,g7670,g12914);
  and AND2_1047(g14007,g7673,g12915);
  and AND2_1048(g14022,g7679,g12921);
  and AND2_1049(g14023,g7682,g12922);
  and AND2_1050(g14039,g7688,g12931);
  and AND2_1051(g14040,g7691,g12932);
  and AND2_1052(g14059,g7697,g12934);
  and AND2_1053(g14067,g7703,g12940);
  and AND2_1054(g14097,g7706,g12943);
  and AND2_1055(g14098,g7709,g12944);
  and AND2_1056(g14113,g7715,g12950);
  and AND2_1057(g14114,g7718,g12951);
  and AND2_1058(g14130,g7724,g12960);
  and AND2_1059(g14131,g7727,g12961);
  and AND2_1060(g14143,g8026,g12965);
  and AND2_1061(g14182,g7733,g12969);
  and AND2_1062(g14212,g7736,g12972);
  and AND2_1063(g14213,g7739,g12973);
  and AND2_1064(g14228,g7745,g12979);
  and AND2_1065(g14229,g7748,g12980);
  and AND2_1066(g14297,g7757,g12993);
  and AND2_1067(g14327,g7760,g12996);
  and AND2_1068(g14328,g7763,g12997);
  and AND2_1069(g14336,g8099,g12998);
  and AND2_1070(g14419,g7779,g13003);
  and AND2_1071(g14690,g7841,g13101);
  and AND2_1072(g14724,g7861,g13117);
  and AND2_1073(g14752,g7891,g13130);
  and AND2_1074(g14767,g13245,g10765);
  and AND2_1075(g14773,g7915,g13141);
  and AND2_1076(g14884,g8169,g12548);
  and AND2_1077(g14894,g3940,g13148);
  and AND2_1078(g14956,g11059,g13151);
  and AND2_1079(g14957,g4015,g13152);
  and AND2_1080(g14958,g4016,g13153);
  and AND2_1081(g14975,g4047,g13154);
  and AND2_1082(g15020,g8090,g12561);
  and AND2_1083(g15030,g4110,g13158);
  and AND2_1084(g15031,g4111,g13159);
  and AND2_1085(g15046,g4142,g13161);
  and AND2_1086(g15047,g4143,g13162);
  and AND2_1087(g15064,g4174,g13163);
  and AND2_1088(g15093,g7869,g12601);
  and AND2_1089(g15094,g7872,g12604);
  and AND2_1090(g15104,g4220,g13167);
  and AND2_1091(g15105,g4224,g13168);
  and AND2_1092(g15126,g4249,g13169);
  and AND2_1093(g15127,g4250,g13170);
  and AND2_1094(g15142,g4281,g13172);
  and AND2_1095(g15143,g4282,g13173);
  and AND2_1096(g15160,g4313,g13174);
  and AND2_1097(g15171,g8015,g12647);
  and AND2_1098(g15172,g4346,g13176);
  and AND2_1099(g15173,g4347,g13177);
  and AND2_1100(g15178,g640,g12651);
  and AND2_1101(g15196,g4375,g13178);
  and AND2_1102(g15197,g4379,g13179);
  and AND2_1103(g15218,g4404,g13180);
  and AND2_1104(g15219,g4405,g13181);
  and AND2_1105(g15234,g4436,g13183);
  and AND2_1106(g15235,g4437,g13184);
  and AND2_1107(g15243,g7849,g12692);
  and AND2_1108(g15244,g7852,g12695);
  and AND2_1109(g15245,g4474,g13185);
  and AND2_1110(g15246,g4475,g13186);
  and AND2_1111(g15247,g4479,g13187);
  and AND2_1112(g15257,g4357,g12702);
  and AND2_1113(g15258,g4515,g13188);
  and AND2_1114(g15259,g4516,g13189);
  and AND2_1115(g15264,g1326,g12705);
  and AND2_1116(g15282,g4544,g13190);
  and AND2_1117(g15283,g4548,g13191);
  and AND2_1118(g15304,g4573,g13192);
  and AND2_1119(g15305,g4574,g13193);
  and AND2_1120(g15320,g7964,g12744);
  and AND2_1121(g15321,g4601,g13195);
  and AND2_1122(g15324,g4609,g13196);
  and AND2_1123(g15325,g4610,g13197);
  and AND2_1124(g15335,g4489,g12749);
  and AND2_1125(g15336,g4492,g12752);
  and AND2_1126(g15337,g4650,g13198);
  and AND2_1127(g15338,g4651,g13199);
  and AND2_1128(g15339,g4655,g13200);
  and AND2_1129(g15349,g4526,g12759);
  and AND2_1130(g15350,g4691,g13201);
  and AND2_1131(g15351,g4692,g13202);
  and AND2_1132(g15356,g2020,g12762);
  and AND2_1133(g15374,g4720,g13203);
  and AND2_1134(g15375,g4724,g13204);
  and AND2_1135(g15388,g7834,g12769);
  and AND2_1136(g15389,g8246,g12772);
  and AND2_1137(g15391,g4752,g13205);
  and AND2_1138(g15392,g4753,g13206);
  and AND2_1139(g15402,g4620,g12783);
  and AND2_1140(g15403,g4623,g12786);
  and AND2_1141(g15407,g4778,g13207);
  and AND2_1142(g15410,g4786,g13208);
  and AND2_1143(g15411,g4787,g13209);
  and AND2_1144(g15421,g4665,g12791);
  and AND2_1145(g15422,g4668,g12794);
  and AND2_1146(g15423,g4827,g13210);
  and AND2_1147(g15424,g4828,g13211);
  and AND2_1148(g15425,g4832,g13212);
  and AND2_1149(g15435,g4702,g12801);
  and AND2_1150(g15436,g4868,g13213);
  and AND2_1151(g15437,g4869,g13214);
  and AND2_1152(g15442,g2714,g12804);
  and AND2_1153(g15452,g7916,g12808);
  and AND2_1154(g15453,g6898,g12811);
  and AND2_1155(g15459,g4897,g13218);
  and AND2_1156(g15460,g4898,g13219);
  and AND2_1157(g15470,g4763,g12816);
  and AND2_1158(g15475,g4928,g13220);
  and AND2_1159(g15476,g4929,g13221);
  and AND2_1160(g15486,g4797,g12822);
  and AND2_1161(g15487,g4800,g12825);
  and AND2_1162(g15491,g4954,g13222);
  and AND2_1163(g15494,g4962,g13223);
  and AND2_1164(g15495,g4963,g13224);
  and AND2_1165(g15505,g4842,g12830);
  and AND2_1166(g15506,g4845,g12833);
  and AND2_1167(g15507,g5003,g13225);
  and AND2_1168(g15508,g5004,g13226);
  and AND2_1169(g15509,g5008,g13227);
  and AND2_1170(g15519,g4879,g12840);
  and AND2_1171(g15520,g8172,g12844);
  and AND2_1172(g15526,g5033,g13232);
  and AND2_1173(g15527,g5034,g13233);
  and AND2_1174(g15545,g5056,g13237);
  and AND2_1175(g15546,g5057,g13238);
  and AND2_1176(g15556,g4939,g12854);
  and AND2_1177(g15561,g5087,g13239);
  and AND2_1178(g15562,g5088,g13240);
  and AND2_1179(g15572,g4973,g12860);
  and AND2_1180(g15573,g4976,g12863);
  and AND2_1181(g15577,g5113,g13241);
  and AND2_1182(g15580,g5121,g13242);
  and AND2_1183(g15581,g5122,g13243);
  and AND2_1184(g15591,g5018,g12868);
  and AND2_1185(g15592,g5021,g12871);
  and AND2_1186(g15593,g7897,g13244);
  and AND2_1187(g15594,g5148,g13249);
  and AND2_1188(g15595,g5149,g13250);
  and AND2_1189(g15604,g5162,g13255);
  and AND2_1190(g15605,g5163,g13256);
  and AND2_1191(g15623,g5185,g13260);
  and AND2_1192(g15624,g5186,g13261);
  and AND2_1193(g15634,g5098,g12895);
  and AND2_1194(g15639,g5216,g13262);
  and AND2_1195(g15640,g5217,g13263);
  and AND2_1196(g15650,g5132,g12901);
  and AND2_1197(g15651,g5135,g12904);
  and AND2_1198(g15658,g8177,g13264);
  and AND2_1199(g15666,g5233,g13268);
  and AND2_1200(g15670,g5241,g13272);
  and AND2_1201(g15671,g5242,g13273);
  and AND2_1202(g15680,g5255,g13278);
  and AND2_1203(g15681,g5256,g13279);
  and AND2_1204(g15699,g5278,g13283);
  and AND2_1205(g15700,g5279,g13284);
  and AND2_1206(g15710,g5227,g12935);
  and AND2_1207(g15717,g7924,g13285);
  and AND2_1208(g15725,g5296,g13293);
  and AND2_1209(g15729,g5304,g13297);
  and AND2_1210(g15730,g5305,g13298);
  and AND2_1211(g15739,g5318,g13303);
  and AND2_1212(g15740,g5319,g13304);
  and AND2_1213(g15753,g7542,g12962);
  and AND2_1214(g15754,g7837,g13308);
  and AND2_1215(g15755,g8178,g13309);
  and AND2_1216(g15765,g5333,g13324);
  and AND2_1217(g15769,g5341,g13328);
  and AND2_1218(g15770,g5342,g13329);
  and AND3_10(II22028,g13004,g3018,g7549);
  and AND3_11(g15780,g7471,g3032,II22028);
  and AND2_1219(g15781,g7971,g13330);
  and AND2_1220(g15793,g5361,g13347);
  and AND2_1221(g15801,g7856,g13351);
  and AND2_1222(g15802,g8253,g13352);
  and AND2_1223(g15817,g8025,g13373);
  and AND2_1224(g15828,g7877,g13398);
  and AND2_1225(g15829,g7857,g13400);
  and AND2_1226(g15840,g8098,g11620);
  and AND2_1227(g15852,g7878,g11642);
  and AND3_12(II22136,g13082,g2912,g7522);
  and AND3_13(g15902,g7607,g2920,II22136);
  and AND2_1228(g15998,g5469,g11732);
  and AND2_1229(g16003,g12013,g10826);
  and AND2_1230(g16004,g5587,g11734);
  and AND2_1231(g16008,g5504,g11735);
  and AND2_1232(g16009,g12071,g10843);
  and AND2_1233(g16010,g7639,g11736);
  and AND2_1234(g16015,g12013,g10859);
  and AND2_1235(g16016,g5601,g11740);
  and AND2_1236(g16017,g12130,g10862);
  and AND2_1237(g16018,g6149,g11741);
  and AND2_1238(g16019,g5507,g11742);
  and AND2_1239(g16028,g5543,g11745);
  and AND2_1240(g16029,g12071,g10877);
  and AND2_1241(g16030,g7667,g11746);
  and AND2_1242(g16031,g6227,g11747);
  and AND2_1243(g16032,g12187,g10883);
  and AND2_1244(g16033,g5546,g11748);
  and AND2_1245(g16045,g12013,g10892);
  and AND2_1246(g16046,g5618,g11761);
  and AND2_1247(g16047,g12130,g10895);
  and AND2_1248(g16048,g6170,g11762);
  and AND2_1249(g16049,g6638,g11763);
  and AND2_1250(g16050,g5590,g11764);
  and AND2_1251(g16051,g12235,g10901);
  and AND2_1252(g16052,g5591,g11765);
  and AND2_1253(g16053,g297,g11770);
  and AND2_1254(g16066,g12071,g10912);
  and AND2_1255(g16067,g7700,g11774);
  and AND2_1256(g16068,g6310,g11775);
  and AND2_1257(g16069,g5346,g11776);
  and AND2_1258(g16070,g12187,g10921);
  and AND2_1259(g16071,g5604,g11777);
  and AND2_1260(g16072,g12275,g10924);
  and AND2_1261(g16073,g5605,g11778);
  and AND2_1262(g16074,g5646,g11782);
  and AND2_1263(g16081,g3304,g11783);
  and AND2_1264(g16089,g984,g11787);
  and AND2_1265(g16100,g12130,g10937);
  and AND2_1266(g16101,g6197,g11794);
  and AND2_1267(g16102,g6905,g11795);
  and AND2_1268(g16103,g5621,g11796);
  and AND2_1269(g16104,g12235,g10946);
  and AND2_1270(g16105,g5622,g11797);
  and AND2_1271(g16106,g12308,g10949);
  and AND2_1272(g16107,g5666,g11801);
  and AND2_1273(g16108,g5667,g11802);
  and AND2_1274(g16109,g8277,g11803);
  and AND2_1275(g16110,g516,g11804);
  and AND2_1276(g16111,g5551,g13215);
  and AND2_1277(g16112,g5684,g11808);
  and AND2_1278(g16119,g3460,g11809);
  and AND2_1279(g16127,g1678,g11813);
  and AND2_1280(g16133,g6444,g11817);
  and AND2_1281(g16134,g5363,g11818);
  and AND2_1282(g16135,g12187,g10980);
  and AND2_1283(g16136,g5640,g11819);
  and AND2_1284(g16137,g12275,g10983);
  and AND2_1285(g16138,g5641,g11820);
  and AND2_1286(g16139,g5704,g11824);
  and AND2_1287(g16140,g5705,g11825);
  and AND2_1288(g16141,g5706,g11826);
  and AND2_1289(g16152,g517,g11829);
  and AND2_1290(g16153,g5592,g13229);
  and AND2_1291(g16158,g5718,g11834);
  and AND2_1292(g16159,g5719,g11835);
  and AND2_1293(g16160,g8286,g11836);
  and AND2_1294(g16161,g1202,g11837);
  and AND2_1295(g16162,g5597,g13234);
  and AND2_1296(g16163,g5736,g11841);
  and AND2_1297(g16170,g3616,g11842);
  and AND2_1298(g16178,g2372,g11846);
  and AND2_1299(g16182,g7149,g11852);
  and AND2_1300(g16183,g12235,g11014);
  and AND2_1301(g16184,g5663,g11853);
  and AND2_1302(g16185,g12308,g11017);
  and AND2_1303(g16186,g5753,g11856);
  and AND2_1304(g16187,g5754,g11857);
  and AND2_1305(g16188,g5755,g11858);
  and AND2_1306(g16197,g518,g11862);
  and AND2_1307(g16198,g5762,g11866);
  and AND2_1308(g16199,g5763,g11867);
  and AND2_1309(g16200,g5764,g11868);
  and AND2_1310(g16211,g1203,g11871);
  and AND2_1311(g16212,g5609,g13252);
  and AND2_1312(g16217,g5776,g11876);
  and AND2_1313(g16218,g5777,g11877);
  and AND2_1314(g16219,g8295,g11878);
  and AND2_1315(g16220,g1896,g11879);
  and AND2_1316(g16221,g5614,g13257);
  and AND2_1317(g16222,g5794,g11883);
  and AND2_1318(g16229,g3772,g11884);
  and AND2_1319(g16237,g5379,g11886);
  and AND2_1320(g16238,g12275,g11066);
  and AND2_1321(g16239,g5700,g11887);
  and AND2_1322(g16240,g5804,g11891);
  and AND2_1323(g16241,g5805,g11892);
  and AND2_1324(g16242,g5806,g11893);
  and AND2_1325(g16250,g519,g11895);
  and AND2_1326(g16251,g5812,g11898);
  and AND2_1327(g16252,g5813,g11899);
  and AND2_1328(g16253,g5814,g11900);
  and AND2_1329(g16262,g1204,g11904);
  and AND2_1330(g16263,g5821,g11908);
  and AND2_1331(g16264,g5822,g11909);
  and AND2_1332(g16265,g5823,g11910);
  and AND2_1333(g16276,g1897,g11913);
  and AND2_1334(g16277,g5634,g13275);
  and AND2_1335(g16282,g5835,g11918);
  and AND2_1336(g16283,g5836,g11919);
  and AND2_1337(g16284,g8304,g11920);
  and AND2_1338(g16285,g2590,g11921);
  and AND2_1339(g16286,g5639,g13280);
  and AND2_1340(g16288,g12308,g11129);
  and AND2_1341(g16289,g5853,g11929);
  and AND2_1342(g16290,g5854,g11930);
  and AND2_1343(g16291,g5855,g11931);
  and AND2_1344(g16292,g294,g11932);
  and AND2_1345(g16298,g520,g11936);
  and AND2_1346(g16299,g5860,g11941);
  and AND2_1347(g16300,g5861,g11942);
  and AND2_1348(g16301,g5862,g11943);
  and AND2_1349(g16309,g1205,g11945);
  and AND2_1350(g16310,g5868,g11948);
  and AND2_1351(g16311,g5869,g11949);
  and AND2_1352(g16312,g5870,g11950);
  and AND2_1353(g16321,g1898,g11954);
  and AND2_1354(g16322,g5877,g11958);
  and AND2_1355(g16323,g5878,g11959);
  and AND2_1356(g16324,g5879,g11960);
  and AND2_1357(g16335,g2591,g11963);
  and AND2_1358(g16336,g5662,g13300);
  and AND2_1359(g16342,g5894,g11968);
  and AND2_1360(g16343,g5895,g11969);
  and AND2_1361(g16344,g5896,g11970);
  and AND2_1362(g16345,g5897,g11971);
  and AND2_1363(g16346,g295,g11972);
  and AND2_1364(g16347,g5900,g11982);
  and AND2_1365(g16348,g5901,g11983);
  and AND2_1366(g16349,g5902,g11984);
  and AND2_1367(g16350,g981,g11985);
  and AND2_1368(g16356,g1206,g11989);
  and AND2_1369(g16357,g5907,g11994);
  and AND2_1370(g16358,g5908,g11995);
  and AND2_1371(g16359,g5909,g11996);
  and AND2_1372(g16367,g1899,g11998);
  and AND2_1373(g16368,g5915,g12001);
  and AND2_1374(g16369,g5916,g12002);
  and AND2_1375(g16370,g5917,g12003);
  and AND2_1376(g16379,g2592,g12007);
  and AND2_1377(g16380,g5925,g12020);
  and AND2_1378(g16381,g5926,g12021);
  and AND2_1379(g16382,g5927,g12022);
  and AND2_1380(g16383,g5928,g12023);
  and AND2_1381(g16384,g296,g12024);
  and AND2_1382(g16385,g5714,g13336);
  and AND2_1383(g16386,g5933,g12037);
  and AND2_1384(g16387,g5934,g12038);
  and AND2_1385(g16388,g5935,g12039);
  and AND2_1386(g16389,g5936,g12040);
  and AND2_1387(g16390,g982,g12041);
  and AND2_1388(g16391,g5939,g12051);
  and AND2_1389(g16392,g5940,g12052);
  and AND2_1390(g16393,g5941,g12053);
  and AND2_1391(g16394,g1675,g12054);
  and AND2_1392(g16400,g1900,g12058);
  and AND2_1393(g16401,g5946,g12063);
  and AND2_1394(g16402,g5947,g12064);
  and AND2_1395(g16403,g5948,g12065);
  and AND2_1396(g16411,g2593,g12067);
  and AND2_1397(g16413,g5954,g12075);
  and AND2_1398(g16414,g5955,g12076);
  and AND2_1399(g16415,g5956,g12077);
  and AND2_1400(g16416,g5957,g12078);
  and AND2_1401(g16417,g5759,g13356);
  and AND2_1402(g16418,g5959,g12084);
  and AND2_1403(g16419,g5960,g12085);
  and AND2_1404(g16420,g5961,g12086);
  and AND2_1405(g16421,g5962,g12087);
  and AND2_1406(g16422,g983,g12088);
  and AND2_1407(g16423,g5772,g13361);
  and AND2_1408(g16424,g5967,g12101);
  and AND2_1409(g16425,g5968,g12102);
  and AND2_1410(g16426,g5969,g12103);
  and AND2_1411(g16427,g5970,g12104);
  and AND2_1412(g16428,g1676,g12105);
  and AND2_1413(g16429,g5973,g12115);
  and AND2_1414(g16430,g5974,g12116);
  and AND2_1415(g16431,g5975,g12117);
  and AND2_1416(g16432,g2369,g12118);
  and AND2_1417(g16438,g2594,g12122);
  and AND2_1418(g16443,g5980,g12134);
  and AND2_1419(g16444,g5981,g12135);
  and AND2_1420(g16445,g5808,g13381);
  and AND2_1421(g16447,g5983,g12147);
  and AND2_1422(g16448,g5984,g12148);
  and AND2_1423(g16449,g5985,g12149);
  and AND2_1424(g16450,g5986,g12150);
  and AND2_1425(g16451,g5818,g13386);
  and AND2_1426(g16452,g5988,g12156);
  and AND2_1427(g16453,g5989,g12157);
  and AND2_1428(g16454,g5990,g12158);
  and AND2_1429(g16455,g5991,g12159);
  and AND2_1430(g16456,g1677,g12160);
  and AND2_1431(g16457,g5831,g13391);
  and AND2_1432(g16458,g5996,g12173);
  and AND2_1433(g16459,g5997,g12174);
  and AND2_1434(g16460,g5998,g12175);
  and AND2_1435(g16461,g5999,g12176);
  and AND2_1436(g16462,g2370,g12177);
  and AND4_22(g16505,g14776,g14797,g16142,g16243);
  and AND4_23(g16513,g15065,g13724,g13764,g13797);
  and AND4_24(g16527,g14811,g14849,g16201,g16302);
  and AND4_25(g16535,g15161,g13774,g13805,g13825);
  and AND4_26(g16558,g14863,g14922,g16266,g16360);
  and AND4_27(g16590,g14936,g15003,g16325,g16404);
  and AND2_1437(g16607,g15022,g15096);
  and AND2_1438(g16625,g15118,g15188);
  and AND2_1439(g16639,g15210,g15274);
  and AND2_1440(g16650,g15296,g15366);
  and AND2_1441(g16850,g6226,g14764);
  and AND2_1442(g16855,g15722,g8646);
  and AND2_1443(g16856,g6443,g14794);
  and AND2_1444(g16859,g15762,g8662);
  and AND2_1445(g16864,g15790,g8681);
  and AND2_1446(g16865,g6896,g14881);
  and AND2_1447(g16879,g15813,g8693);
  and AND2_1448(g16894,g7156,g14959);
  and AND2_1449(g16907,g7335,g15017);
  and AND2_1450(g16908,g7838,g15032);
  and AND2_1451(g16909,g6908,g15033);
  and AND2_1452(g16923,g7352,g15048);
  and AND2_1453(g16938,g7858,g15128);
  and AND2_1454(g16939,g7158,g15129);
  and AND2_1455(g16953,g7482,g15144);
  and AND2_1456(g16964,g7520,g15170);
  and AND2_1457(g16966,g7529,g15174);
  and AND2_1458(g16967,g7827,g15175);
  and AND2_1459(g16968,g6672,g15176);
  and AND2_1460(g16969,g7888,g15220);
  and AND2_1461(g16970,g7354,g15221);
  and AND2_1462(g16984,g7538,g15236);
  and AND2_1463(g16987,g7555,g15260);
  and AND2_1464(g16988,g7842,g15261);
  and AND2_1465(g16989,g6974,g15262);
  and AND2_1466(g16990,g7912,g15306);
  and AND2_1467(g16991,g7484,g15307);
  and AND2_1468(g16993,g7576,g15322);
  and AND2_1469(g16994,g7819,g15323);
  and AND2_1470(g16997,g7578,g15352);
  and AND2_1471(g16998,g7862,g15353);
  and AND2_1472(g16999,g7224,g15354);
  and AND3_14(g17001,g3254,g10694,g14144);
  and AND2_1473(g17015,g7996,g15390);
  and AND2_1474(g17017,g7590,g15408);
  and AND2_1475(g17018,g7830,g15409);
  and AND2_1476(g17021,g7592,g15438);
  and AND2_1477(g17022,g7892,g15439);
  and AND2_1478(g17023,g7420,g15440);
  and AND2_1479(g17028,g7604,g15458);
  and AND3_15(g17031,g3410,g10714,g14259);
  and AND2_1480(g17045,g8071,g15474);
  and AND2_1481(g17047,g7605,g15492);
  and AND2_1482(g17048,g7845,g15493);
  and AND2_1483(g17055,g7153,g15524);
  and AND2_1484(g17056,g7953,g15525);
  and AND2_1485(g17062,g7613,g15544);
  and AND3_16(g17065,g3566,g10735,g14381);
  and AND2_1486(g17079,g8156,g15560);
  and AND2_1487(g17081,g7614,g15578);
  and AND2_1488(g17082,g7865,g15579);
  and AND2_1489(g17084,g7629,g13954);
  and AND2_1490(g17090,g7349,g15602);
  and AND2_1491(g17091,g8004,g15603);
  and AND2_1492(g17097,g7622,g15622);
  and AND3_17(g17100,g3722,g10754,g14493);
  and AND2_1493(g17114,g8242,g15638);
  and AND2_1494(g17116,g7649,g14008);
  and AND2_1495(g17117,g7906,g15665);
  and AND2_1496(g17122,g7658,g14024);
  and AND2_1497(g17128,g7479,g15678);
  and AND2_1498(g17129,g8079,g15679);
  and AND2_1499(g17135,g7638,g15698);
  and AND2_1500(g17138,g7676,g14068);
  and AND2_1501(g17143,g7685,g14099);
  and AND2_1502(g17144,g7958,g15724);
  and AND2_1503(g17149,g7694,g14115);
  and AND2_1504(g17155,g7535,g15737);
  and AND2_1505(g17156,g8164,g15738);
  and AND2_1506(g17161,g7712,g14183);
  and AND2_1507(g17166,g7721,g14214);
  and AND2_1508(g17167,g8009,g15764);
  and AND2_1509(g17172,g7730,g14230);
  and AND2_1510(g17176,g7742,g14298);
  and AND2_1511(g17181,g7751,g14329);
  and AND2_1512(g17182,g8084,g15792);
  and AND2_1513(g17193,g7766,g14420);
  and AND2_1514(g17268,g8024,g15991);
  and AND2_1515(g17301,g8097,g15994);
  and AND2_1516(g17339,g8176,g15997);
  and AND2_1517(g17352,g3942,g14960);
  and AND2_1518(g17353,g3945,g14963);
  and AND2_1519(g17381,g8250,g16001);
  and AND2_1520(g17382,g8252,g16002);
  and AND2_1521(g17393,g3941,g16005);
  and AND2_1522(g17395,g6177,g15034);
  and AND2_1523(g17396,g4020,g15037);
  and AND2_1524(g17397,g4023,g15040);
  and AND2_1525(g17398,g4026,g15043);
  and AND2_1526(g17408,g4049,g15049);
  and AND2_1527(g17409,g4052,g15052);
  and AND2_1528(g17428,g3994,g16007);
  and AND2_1529(g17446,g6284,g16011);
  and AND2_1530(g17447,g4115,g15106);
  and AND2_1531(g17448,g4118,g15109);
  and AND2_1532(g17449,g4121,g15112);
  and AND2_1533(g17450,g4124,g15115);
  and AND2_1534(g17460,g4048,g16012);
  and AND2_1535(g17461,g6209,g15130);
  and AND2_1536(g17462,g4147,g15133);
  and AND2_1537(g17463,g4150,g15136);
  and AND2_1538(g17464,g4153,g15139);
  and AND2_1539(g17474,g4176,g15145);
  and AND2_1540(g17475,g4179,g15148);
  and AND2_1541(g17485,g4089,g16013);
  and AND2_1542(g17486,g4091,g16014);
  and AND2_1543(g17506,g6675,g16023);
  and AND2_1544(g17508,g4225,g15179);
  and AND2_1545(g17509,g4228,g15182);
  and AND2_1546(g17510,g4231,g15185);
  and AND2_1547(g17526,g6421,g16025);
  and AND2_1548(g17527,g4254,g15198);
  and AND2_1549(g17528,g4257,g15201);
  and AND2_1550(g17529,g4260,g15204);
  and AND2_1551(g17530,g4263,g15207);
  and AND2_1552(g17540,g4175,g16026);
  and AND2_1553(g17541,g6298,g15222);
  and AND2_1554(g17542,g4286,g15225);
  and AND2_1555(g17543,g4289,g15228);
  and AND2_1556(g17544,g4292,g15231);
  and AND2_1557(g17554,g4315,g15237);
  and AND2_1558(g17555,g4318,g15240);
  and AND2_1559(g17556,g4201,g16027);
  and AND2_1560(g17576,g4348,g15248);
  and AND2_1561(g17577,g4351,g15251);
  and AND2_1562(g17578,g4354,g15254);
  and AND2_1563(g17597,g6977,g16039);
  and AND2_1564(g17598,g4380,g15265);
  and AND2_1565(g17599,g4383,g15268);
  and AND2_1566(g17600,g4386,g15271);
  and AND2_1567(g17616,g6626,g16041);
  and AND2_1568(g17617,g4409,g15284);
  and AND2_1569(g17618,g4412,g15287);
  and AND2_1570(g17619,g4415,g15290);
  and AND2_1571(g17620,g4418,g15293);
  and AND2_1572(g17630,g4314,g16042);
  and AND2_1573(g17631,g6435,g15308);
  and AND2_1574(g17632,g4441,g15311);
  and AND2_1575(g17633,g4444,g15314);
  and AND2_1576(g17634,g4447,g15317);
  and AND2_1577(g17635,g4322,g16043);
  and AND2_1578(g17636,g4324,g16044);
  and AND2_1579(g17652,g4480,g15326);
  and AND2_1580(g17653,g4483,g15329);
  and AND2_1581(g17654,g4486,g15332);
  and AND2_1582(g17673,g4517,g15340);
  and AND2_1583(g17674,g4520,g15343);
  and AND2_1584(g17675,g4523,g15346);
  and AND2_1585(g17694,g7227,g16061);
  and AND2_1586(g17695,g4549,g15357);
  and AND2_1587(g17696,g4552,g15360);
  and AND2_1588(g17697,g4555,g15363);
  and AND2_1589(g17713,g6890,g16063);
  and AND2_1590(g17714,g4578,g15376);
  and AND2_1591(g17715,g4581,g15379);
  and AND2_1592(g17716,g4584,g15382);
  and AND2_1593(g17717,g4587,g15385);
  and AND2_1594(g17718,g4451,g16064);
  and AND2_1595(g17719,g2993,g16065);
  and AND2_1596(g17734,g4611,g15393);
  and AND2_1597(g17735,g4614,g15396);
  and AND2_1598(g17736,g4617,g15399);
  and AND2_1599(g17737,g4626,g15404);
  and AND2_1600(g17752,g4656,g15412);
  and AND2_1601(g17753,g4659,g15415);
  and AND2_1602(g17754,g4662,g15418);
  and AND2_1603(g17773,g4693,g15426);
  and AND2_1604(g17774,g4696,g15429);
  and AND2_1605(g17775,g4699,g15432);
  and AND2_1606(g17794,g7423,g16097);
  and AND2_1607(g17795,g4725,g15443);
  and AND2_1608(g17796,g4728,g15446);
  and AND2_1609(g17797,g4731,g15449);
  and AND2_1610(g17798,g4591,g16099);
  and AND2_1611(g17812,g4754,g15461);
  and AND2_1612(g17813,g4757,g15464);
  and AND2_1613(g17814,g4760,g15467);
  and AND2_1614(g17824,g4766,g15471);
  and AND2_1615(g17835,g4788,g15477);
  and AND2_1616(g17836,g4791,g15480);
  and AND2_1617(g17837,g4794,g15483);
  and AND2_1618(g17838,g4803,g15488);
  and AND2_1619(g17853,g4833,g15496);
  and AND2_1620(g17854,g4836,g15499);
  and AND2_1621(g17855,g4839,g15502);
  and AND2_1622(g17874,g4870,g15510);
  and AND2_1623(g17875,g4873,g15513);
  and AND2_1624(g17876,g4876,g15516);
  and AND2_1625(g17877,g2998,g15521);
  and AND2_1626(g17900,g4899,g15528);
  and AND2_1627(g17901,g4902,g15531);
  and AND2_1628(g17902,g4905,g15534);
  and AND2_1629(g17912,g4908,g15537);
  and AND2_1630(g17924,g4930,g15547);
  and AND2_1631(g17925,g4933,g15550);
  and AND2_1632(g17926,g4936,g15553);
  and AND2_1633(g17936,g4942,g15557);
  and AND2_1634(g17947,g4964,g15563);
  and AND2_1635(g17948,g4967,g15566);
  and AND2_1636(g17949,g4970,g15569);
  and AND2_1637(g17950,g4979,g15574);
  and AND2_1638(g17965,g5009,g15582);
  and AND2_1639(g17966,g5012,g15585);
  and AND2_1640(g17967,g5015,g15588);
  and AND2_1641(g17989,g5035,g15596);
  and AND2_1642(g17990,g5038,g15599);
  and AND2_1643(g18011,g5058,g15606);
  and AND2_1644(g18012,g5061,g15609);
  and AND2_1645(g18013,g5064,g15612);
  and AND2_1646(g18023,g5067,g15615);
  and AND2_1647(g18035,g5089,g15625);
  and AND2_1648(g18036,g5092,g15628);
  and AND2_1649(g18037,g5095,g15631);
  and AND2_1650(g18047,g5101,g15635);
  and AND2_1651(g18058,g5123,g15641);
  and AND2_1652(g18059,g5126,g15644);
  and AND2_1653(g18060,g5129,g15647);
  and AND2_1654(g18061,g5138,g15652);
  and AND2_1655(g18062,g7462,g15655);
  and AND2_1656(g18088,g5150,g15667);
  and AND2_1657(g18106,g5164,g15672);
  and AND2_1658(g18107,g5167,g15675);
  and AND2_1659(g18128,g5187,g15682);
  and AND2_1660(g18129,g5190,g15685);
  and AND2_1661(g18130,g5193,g15688);
  and AND2_1662(g18140,g5196,g15691);
  and AND2_1663(g18152,g5218,g15701);
  and AND2_1664(g18153,g5221,g15704);
  and AND2_1665(g18154,g5224,g15707);
  and AND2_1666(g18164,g5230,g15711);
  and AND2_1667(g18165,g2883,g16287);
  and AND2_1668(g18169,g7527,g15714);
  and AND2_1669(g18204,g5243,g15726);
  and AND2_1670(g18222,g5257,g15731);
  and AND2_1671(g18223,g5260,g15734);
  and AND2_1672(g18244,g5280,g15741);
  and AND2_1673(g18245,g5283,g15744);
  and AND2_1674(g18246,g5286,g15747);
  and AND2_1675(g18256,g5289,g15750);
  and AND2_1676(g18311,g5306,g15766);
  and AND2_1677(g18329,g5320,g15771);
  and AND2_1678(g18330,g5323,g15774);
  and AND2_1679(g18333,g2888,g15777);
  and AND2_1680(g18404,g5343,g15794);
  and AND3_18(II24619,g14776,g14837,g16142);
  and AND3_19(g18547,g13677,g13750,II24619);
  and AND3_20(II24689,g14811,g14910,g16201);
  and AND3_21(g18597,g13714,g13791,II24689);
  and AND3_22(II24738,g14863,g14991,g16266);
  and AND3_23(g18629,g13764,g13819,II24738);
  and AND3_24(II24758,g14936,g15080,g16325);
  and AND3_25(g18638,g13805,g13840,II24758);
  and AND4_28(g18645,g14776,g14895,g16142,g13750);
  and AND3_26(g18647,g14895,g16142,g16243);
  and AND4_29(g18648,g14811,g14976,g16201,g13791);
  and AND4_30(g18649,g14776,g14837,g13657,g16189);
  and AND3_27(g18650,g14976,g16201,g16302);
  and AND4_31(g18651,g14863,g15065,g16266,g13819);
  and AND4_32(g18652,g14797,g13657,g13677,g16243);
  and AND4_33(g18653,g14811,g14910,g13687,g16254);
  and AND3_28(g18654,g15065,g16266,g16360);
  and AND4_34(g18655,g14936,g15161,g16325,g13840);
  and AND4_35(g18665,g14776,g14837,g16189,g13706);
  and AND4_36(g18666,g14849,g13687,g13714,g16302);
  and AND4_37(g18667,g14863,g14991,g13724,g16313);
  and AND3_29(g18668,g15161,g16325,g16404);
  and AND4_38(g18688,g14811,g14910,g16254,g13756);
  and AND4_39(g18689,g14922,g13724,g13764,g16360);
  and AND4_40(g18690,g14936,g15080,g13774,g16371);
  and AND4_41(g18717,g14863,g14991,g16313,g13797);
  and AND4_42(g18718,g15003,g13774,g13805,g16404);
  and AND4_43(g18753,g14936,g15080,g16371,g13825);
  and AND2_1681(g18982,g13519,g16154);
  and AND2_1682(g18990,g13530,g16213);
  and AND4_44(g18994,g14895,g13657,g13677,g13706);
  and AND2_1683(g18997,g13541,g16278);
  and AND4_45(g19007,g14976,g13687,g13714,g13756);
  and AND2_1684(g19010,g13552,g16337);
  and AND4_46(g19063,g18679,g14910,g13687,g16254);
  and AND4_47(g19079,g14797,g18692,g16142,g16189);
  and AND4_48(g19080,g18708,g14991,g13724,g16313);
  and AND2_1685(g19087,g17215,g16540);
  and AND4_49(g19088,g18656,g14797,g16189,g13706);
  and AND4_50(g19089,g14849,g18728,g16201,g16254);
  and AND4_51(g19090,g18744,g15080,g13774,g16371);
  and AND4_52(g19092,g14776,g18670,g18692,g16293);
  and AND2_1686(g19093,g17218,g16572);
  and AND4_53(g19094,g18679,g14849,g16254,g13756);
  and AND4_54(g19095,g14922,g18765,g16266,g16313);
  and AND3_30(II25280,g18656,g18670,g18720);
  and AND3_31(g19097,g13657,g16243,II25280);
  and AND4_55(g19099,g14811,g18699,g18728,g16351);
  and AND2_1687(g19100,g17220,g16596);
  and AND4_56(g19101,g18708,g14922,g16313,g13797);
  and AND4_57(g19102,g15003,g18796,g16325,g16371);
  and AND3_32(II25291,g18679,g18699,g18758);
  and AND3_33(g19104,g13687,g16302,II25291);
  and AND4_58(g19106,g14863,g18735,g18765,g16395);
  and AND2_1688(g19107,g17223,g16616);
  and AND4_59(g19108,g18744,g15003,g16371,g13825);
  and AND3_34(II25300,g18708,g18735,g18789);
  and AND3_35(g19109,g13724,g16360,II25300);
  and AND4_60(g19111,g14936,g18772,g18796,g16433);
  and AND2_1689(g19112,g14657,g16633);
  and AND3_36(II25311,g18744,g18772,g18815);
  and AND3_37(g19116,g13774,g16404,II25311);
  and AND2_1690(g19117,g14691,g16644);
  and AND2_1691(g19124,g14725,g16656);
  and AND2_1692(g19131,g14753,g16673);
  and AND2_1693(g19142,g17159,g16719);
  and AND2_1694(g19143,g17174,g16761);
  and AND2_1695(g19146,g17191,g16788);
  and AND2_1696(g19148,g17202,g16817);
  and AND2_1697(g19150,g17189,g8602);
  and AND2_1698(g19155,g17200,g8614);
  and AND2_1699(g19161,g17207,g8627);
  and AND2_1700(g19166,g17212,g8637);
  and AND2_1701(g19228,g16662,g12125);
  and AND2_1702(g19236,g16935,g8802);
  and AND3_38(g19241,g16867,g14158,g14071);
  and AND2_1703(g19248,g16662,g8817);
  and AND2_1704(g19252,g18725,g9527);
  and AND3_39(g19254,g16895,g14273,g14186);
  and AND2_1705(g19260,g16749,g3124);
  and AND3_40(g19267,g16924,g14395,g14301);
  and AND3_41(g19282,g16954,g14507,g14423);
  and AND2_1706(g19284,g18063,g3111);
  and AND2_1707(g19285,g16749,g7642);
  and AND2_1708(g19289,g17029,g8580);
  and AND3_42(g19303,g16867,g16543,g14071);
  and AND2_1709(g19307,g17063,g8587);
  and AND2_1710(g19316,g18063,g3110);
  and AND2_1711(g19317,g16749,g3126);
  and AND3_43(g19320,g16867,g16515,g14158);
  and AND3_44(g19324,g16895,g16575,g14186);
  and AND2_1712(g19328,g17098,g8594);
  and AND3_45(g19347,g16895,g16546,g14273);
  and AND3_46(g19351,g16924,g16599,g14301);
  and AND2_1713(g19355,g17136,g8605);
  and AND2_1714(g19356,g18063,g3112);
  and AND3_47(g19381,g16924,g16578,g14395);
  and AND3_48(g19385,g16954,g16619,g14423);
  and AND3_49(g19413,g16954,g16602,g14507);
  and AND3_50(g19449,g16884,g14797,g14776);
  and AND3_51(g19476,g16913,g14849,g14811);
  and AND3_52(g19499,g16943,g14922,g14863);
  and AND3_53(g19520,g16974,g15003,g14936);
  and AND3_54(g19531,g16884,g16722,g14776);
  and AND3_55(g19540,g16884,g16697,g14797);
  and AND3_56(g19541,g16913,g16764,g14811);
  and AND3_57(g19544,g16913,g16728,g14849);
  and AND3_58(g19545,g16943,g16791,g14863);
  and AND3_59(g19547,g16943,g16770,g14922);
  and AND3_60(g19548,g16974,g16820,g14936);
  and AND2_1715(g19549,g7950,g17230);
  and AND3_61(g19551,g16974,g16797,g15003);
  and AND2_1716(g19552,g16829,g6048);
  and AND2_1717(g19553,g7990,g17237);
  and AND2_1718(g19554,g7993,g17240);
  and AND2_1719(g19555,g8001,g17243);
  and AND2_1720(g19557,g8053,g17249);
  and AND2_1721(g19558,g8056,g17252);
  and AND2_1722(g19559,g8059,g17255);
  and AND2_1723(g19560,g8065,g17259);
  and AND2_1724(g19561,g8068,g17262);
  and AND2_1725(g19562,g8076,g17265);
  and AND2_1726(g19564,g8123,g17272);
  and AND2_1727(g19565,g8126,g17275);
  and AND2_1728(g19566,g8129,g17278);
  and AND2_1729(g19567,g8138,g17282);
  and AND2_1730(g19568,g8141,g17285);
  and AND2_1731(g19569,g8144,g17288);
  and AND2_1732(g19570,g8150,g17291);
  and AND2_1733(g19571,g8153,g17294);
  and AND2_1734(g19572,g8161,g17297);
  and AND2_1735(g19574,g8191,g17304);
  and AND2_1736(g19575,g8194,g17307);
  and AND2_1737(g19576,g8197,g17310);
  and AND2_1738(g19584,g640,g18756);
  and AND2_1739(g19585,g692,g18757);
  and AND2_1740(g19586,g8209,g17315);
  and AND2_1741(g19587,g8212,g17318);
  and AND2_1742(g19588,g8215,g17321);
  and AND2_1743(g19589,g8224,g17324);
  and AND2_1744(g19590,g8227,g17327);
  and AND2_1745(g19591,g8230,g17330);
  and AND2_1746(g19592,g8236,g17333);
  and AND2_1747(g19593,g8239,g17336);
  and AND2_1748(g19594,g16935,g12555);
  and AND2_1749(g19597,g3922,g17342);
  and AND2_1750(g19598,g3925,g17345);
  and AND2_1751(g19599,g3928,g17348);
  and AND2_1752(g19600,g633,g18783);
  and AND2_1753(g19601,g640,g18784);
  and AND2_1754(g19602,g633,g18785);
  and AND2_1755(g19603,g692,g18786);
  and AND2_1756(g19604,g3948,g17354);
  and AND2_1757(g19605,g3951,g17357);
  and AND2_1758(g19606,g3954,g17360);
  and AND2_1759(g19614,g1326,g18787);
  and AND2_1760(g19615,g1378,g18788);
  and AND2_1761(g19616,g3966,g17363);
  and AND2_1762(g19617,g3969,g17366);
  and AND2_1763(g19618,g3972,g17369);
  and AND2_1764(g19619,g3981,g17372);
  and AND2_1765(g19620,g3984,g17375);
  and AND2_1766(g19621,g3987,g17378);
  and AND2_1767(g19623,g4000,g17384);
  and AND2_1768(g19624,g4003,g17387);
  and AND2_1769(g19625,g4006,g17390);
  and AND2_1770(g19626,g640,g18805);
  and AND2_1771(g19627,g633,g18806);
  and AND2_1772(g19628,g653,g18807);
  and AND2_1773(g19629,g692,g18808);
  and AND2_1774(g19630,g4029,g17399);
  and AND2_1775(g19631,g4032,g17402);
  and AND2_1776(g19632,g4035,g17405);
  and AND2_1777(g19633,g1319,g18809);
  and AND2_1778(g19634,g1326,g18810);
  and AND2_1779(g19635,g1319,g18811);
  and AND2_1780(g19636,g1378,g18812);
  and AND2_1781(g19637,g4055,g17410);
  and AND2_1782(g19638,g4058,g17413);
  and AND2_1783(g19639,g4061,g17416);
  and AND2_1784(g19647,g2020,g18813);
  and AND2_1785(g19648,g2072,g18814);
  and AND2_1786(g19649,g4073,g17419);
  and AND2_1787(g19650,g4076,g17422);
  and AND2_1788(g19651,g4079,g17425);
  and AND2_1789(g19653,g4095,g17430);
  and AND2_1790(g19654,g4098,g17433);
  and AND2_1791(g19655,g4101,g17436);
  and AND2_1792(g19656,g4104,g17439);
  and AND2_1793(g19660,g633,g18822);
  and AND2_1794(g19661,g653,g18823);
  and AND2_1795(g19662,g646,g18824);
  and AND2_1796(g19663,g4127,g17451);
  and AND2_1797(g19664,g4130,g17454);
  and AND2_1798(g19665,g4133,g17457);
  and AND2_1799(g19666,g1326,g18825);
  and AND2_1800(g19667,g1319,g18826);
  and AND2_1801(g19668,g1339,g18827);
  and AND2_1802(g19669,g1378,g18828);
  and AND2_1803(g19670,g4156,g17465);
  and AND2_1804(g19671,g4159,g17468);
  and AND2_1805(g19672,g4162,g17471);
  and AND2_1806(g19673,g2013,g18829);
  and AND2_1807(g19674,g2020,g18830);
  and AND2_1808(g19675,g2013,g18831);
  and AND2_1809(g19676,g2072,g18832);
  and AND2_1810(g19677,g4182,g17476);
  and AND2_1811(g19678,g4185,g17479);
  and AND2_1812(g19679,g4188,g17482);
  and AND2_1813(g19687,g2714,g18833);
  and AND2_1814(g19688,g2766,g18834);
  and AND2_1815(g19691,g16841,g10865);
  and AND2_1816(g19692,g4205,g17487);
  and AND2_1817(g19693,g4208,g17490);
  and AND2_1818(g19694,g4211,g17493);
  and AND2_1819(g19695,g4214,g17496);
  and AND2_1820(g19697,g653,g18838);
  and AND2_1821(g19698,g646,g18839);
  and AND2_1822(g19699,g660,g18840);
  and AND2_1823(g19700,g17815,g16024);
  and AND2_1824(g19701,g4234,g17511);
  and AND2_1825(g19702,g4237,g17514);
  and AND2_1826(g19703,g4240,g17517);
  and AND2_1827(g19704,g4243,g17520);
  and AND2_1828(g19708,g1319,g18841);
  and AND2_1829(g19709,g1339,g18842);
  and AND2_1830(g19710,g1332,g18843);
  and AND2_1831(g19711,g4266,g17531);
  and AND2_1832(g19712,g4269,g17534);
  and AND2_1833(g19713,g4272,g17537);
  and AND2_1834(g19714,g2020,g18844);
  and AND2_1835(g19715,g2013,g18845);
  and AND2_1836(g19716,g2033,g18846);
  and AND2_1837(g19717,g2072,g18847);
  and AND2_1838(g19718,g4295,g17545);
  and AND2_1839(g19719,g4298,g17548);
  and AND2_1840(g19720,g4301,g17551);
  and AND2_1841(g19721,g2707,g18848);
  and AND2_1842(g19722,g2714,g18849);
  and AND2_1843(g19723,g2707,g18850);
  and AND2_1844(g19724,g2766,g18851);
  and AND2_1845(g19726,g16847,g6131);
  and AND2_1846(g19727,g4329,g17557);
  and AND2_1847(g19728,g4332,g17560);
  and AND2_1848(g19729,g4335,g17563);
  and AND2_1849(g19730,g653,g17573);
  and AND2_1850(g19731,g646,g18853);
  and AND2_1851(g19732,g660,g18854);
  and AND2_1852(g19733,g672,g18855);
  and AND2_1853(g19734,g17815,g16034);
  and AND2_1854(g19735,g17903,g16035);
  and AND2_1855(g19736,g4360,g17579);
  and AND2_1856(g19737,g4363,g17582);
  and AND2_1857(g19738,g4366,g17585);
  and AND2_1858(g19739,g4369,g17588);
  and AND2_1859(g19741,g1339,g18856);
  and AND2_1860(g19742,g1332,g18857);
  and AND2_1861(g19743,g1346,g18858);
  and AND2_1862(g19744,g17927,g16040);
  and AND2_1863(g19745,g4389,g17601);
  and AND2_1864(g19746,g4392,g17604);
  and AND2_1865(g19747,g4395,g17607);
  and AND2_1866(g19748,g4398,g17610);
  and AND2_1867(g19752,g2013,g18859);
  and AND2_1868(g19753,g2033,g18860);
  and AND2_1869(g19754,g2026,g18861);
  and AND2_1870(g19755,g4421,g17621);
  and AND2_1871(g19756,g4424,g17624);
  and AND2_1872(g19757,g4427,g17627);
  and AND2_1873(g19758,g2714,g18862);
  and AND2_1874(g19759,g2707,g18863);
  and AND2_1875(g19760,g2727,g18864);
  and AND2_1876(g19761,g2766,g18865);
  and AND2_1877(g19764,g4453,g17637);
  and AND2_1878(g19765,g660,g18870);
  and AND2_1879(g19766,g672,g18871);
  and AND2_1880(g19767,g666,g18872);
  and AND2_1881(g19768,g17815,g16054);
  and AND2_1882(g19769,g17903,g16055);
  and AND2_1883(g19770,g4498,g17655);
  and AND2_1884(g19771,g4501,g17658);
  and AND2_1885(g19772,g4504,g17661);
  and AND2_1886(g19773,g1339,g17670);
  and AND2_1887(g19774,g1332,g18874);
  and AND2_1888(g19775,g1346,g18875);
  and AND2_1889(g19776,g1358,g18876);
  and AND2_1890(g19777,g17927,g16056);
  and AND2_1891(g19778,g18014,g16057);
  and AND2_1892(g19779,g4529,g17676);
  and AND2_1893(g19780,g4532,g17679);
  and AND2_1894(g19781,g4535,g17682);
  and AND2_1895(g19782,g4538,g17685);
  and AND2_1896(g19784,g2033,g18877);
  and AND2_1897(g19785,g2026,g18878);
  and AND2_1898(g19786,g2040,g18879);
  and AND2_1899(g19787,g18038,g16062);
  and AND2_1900(g19788,g4558,g17698);
  and AND2_1901(g19789,g4561,g17701);
  and AND2_1902(g19790,g4564,g17704);
  and AND2_1903(g19791,g4567,g17707);
  and AND2_1904(g19795,g2707,g18880);
  and AND2_1905(g19796,g2727,g18881);
  and AND2_1906(g19797,g2720,g18882);
  and AND3_62(II26240,g18174,g18341,g17974);
  and AND3_63(g19799,g17640,g18074,II26240);
  and AND2_1907(g19802,g672,g18891);
  and AND2_1908(g19803,g666,g18892);
  and AND2_1909(g19804,g679,g18893);
  and AND2_1910(g19805,g17903,g16088);
  and AND2_1911(g19806,g4629,g17738);
  and AND2_1912(g19807,g1346,g18896);
  and AND2_1913(g19808,g1358,g18897);
  and AND2_1914(g19809,g1352,g18898);
  and AND2_1915(g19810,g17927,g16090);
  and AND2_1916(g19811,g18014,g16091);
  and AND2_1917(g19812,g4674,g17755);
  and AND2_1918(g19813,g4677,g17758);
  and AND2_1919(g19814,g4680,g17761);
  and AND2_1920(g19815,g2033,g17770);
  and AND2_1921(g19816,g2026,g18900);
  and AND2_1922(g19817,g2040,g18901);
  and AND2_1923(g19818,g2052,g18902);
  and AND2_1924(g19819,g18038,g16092);
  and AND2_1925(g19820,g18131,g16093);
  and AND2_1926(g19821,g4705,g17776);
  and AND2_1927(g19822,g4708,g17779);
  and AND2_1928(g19823,g4711,g17782);
  and AND2_1929(g19824,g4714,g17785);
  and AND2_1930(g19826,g2727,g18903);
  and AND2_1931(g19827,g2720,g18904);
  and AND2_1932(g19828,g2734,g18905);
  and AND2_1933(g19829,g18155,g16098);
  and AND2_1934(g19836,g7143,g18908);
  and AND2_1935(g19837,g6901,g17799);
  and AND2_1936(g19839,g666,g18909);
  and AND2_1937(g19840,g679,g18910);
  and AND2_1938(g19841,g686,g18911);
  and AND3_64(II26282,g18188,g18089,g17991);
  and AND3_65(g19842,g14525,g13922,II26282);
  and AND3_66(II26285,g18281,g18436,g18091);
  and AND3_67(g19843,g17741,g18190,II26285);
  and AND2_1939(g19846,g1358,g18914);
  and AND2_1940(g19847,g1352,g18915);
  and AND2_1941(g19848,g1365,g18916);
  and AND2_1942(g19849,g18014,g16126);
  and AND2_1943(g19850,g4806,g17839);
  and AND2_1944(g19851,g2040,g18919);
  and AND2_1945(g19852,g2052,g18920);
  and AND2_1946(g19853,g2046,g18921);
  and AND2_1947(g19854,g18038,g16128);
  and AND2_1948(g19855,g18131,g16129);
  and AND2_1949(g19856,g4851,g17856);
  and AND2_1950(g19857,g4854,g17859);
  and AND2_1951(g19858,g4857,g17862);
  and AND2_1952(g19859,g2727,g17871);
  and AND2_1953(g19860,g2720,g18923);
  and AND2_1954(g19861,g2734,g18924);
  and AND2_1955(g19862,g2746,g18925);
  and AND2_1956(g19863,g18155,g16130);
  and AND2_1957(g19864,g18247,g16131);
  and AND3_68(g19868,g16498,g16867,g19001);
  and AND2_1958(g19869,g679,g18926);
  and AND2_1959(g19870,g686,g18927);
  and AND3_69(II26311,g18353,g13958,g14011);
  and AND3_70(g19871,g14086,g18275,II26311);
  and AND2_1960(g19872,g1352,g18928);
  and AND2_1961(g19873,g1365,g18929);
  and AND2_1962(g19874,g1372,g18930);
  and AND3_71(II26317,g18295,g18205,g18108);
  and AND3_72(g19875,g14580,g13978,II26317);
  and AND3_73(II26320,g18374,g18509,g18207);
  and AND3_74(g19876,g17842,g18297,II26320);
  and AND2_1963(g19879,g2052,g18933);
  and AND2_1964(g19880,g2046,g18934);
  and AND2_1965(g19881,g2059,g18935);
  and AND2_1966(g19882,g18131,g16177);
  and AND2_1967(g19883,g4982,g17951);
  and AND2_1968(g19884,g2734,g18938);
  and AND2_1969(g19885,g2746,g18939);
  and AND2_1970(g19886,g2740,g18940);
  and AND2_1971(g19887,g18155,g16179);
  and AND2_1972(g19888,g18247,g16180);
  and AND2_1973(g19889,g2912,g18943);
  and AND2_1974(g19895,g686,g18945);
  and AND3_75(g19899,g16520,g16895,g16507);
  and AND2_1975(g19900,g1365,g18946);
  and AND2_1976(g19901,g1372,g18947);
  and AND3_76(II26348,g18448,g14028,g14102);
  and AND3_77(g19902,g14201,g18368,II26348);
  and AND2_1977(g19903,g2046,g18948);
  and AND2_1978(g19904,g2059,g18949);
  and AND2_1979(g19905,g2066,g18950);
  and AND3_78(II26354,g18388,g18312,g18224);
  and AND3_79(g19906,g14614,g14048,II26354);
  and AND3_80(II26357,g18469,g18573,g18314);
  and AND3_81(g19907,g17954,g18390,II26357);
  and AND2_1980(g19910,g2746,g18953);
  and AND2_1981(g19911,g2740,g18954);
  and AND2_1982(g19912,g2753,g18955);
  and AND2_1983(g19913,g18247,g16236);
  and AND2_1984(g19914,g3018,g18958);
  and AND2_1985(g19920,g1372,g18961);
  and AND3_82(g19924,g16551,g16924,g16529);
  and AND2_1986(g19925,g2059,g18962);
  and AND2_1987(g19926,g2066,g18963);
  and AND3_83(II26377,g18521,g14119,g14217);
  and AND3_84(g19927,g14316,g18463,II26377);
  and AND2_1988(g19928,g2740,g18964);
  and AND2_1989(g19929,g2753,g18965);
  and AND2_1990(g19930,g2760,g18966);
  and AND3_85(II26383,g18483,g18405,g18331);
  and AND3_86(g19931,g14637,g14139,II26383);
  and AND2_1991(g19932,g2917,g18166);
  and AND2_1992(g19935,g2066,g18972);
  and AND3_87(g19939,g16583,g16954,g16560);
  and AND2_1993(g19940,g2753,g18973);
  and AND2_1994(g19941,g2760,g18974);
  and AND3_88(II26396,g18585,g14234,g14332);
  and AND3_89(g19942,g14438,g18536,II26396);
  and AND2_1995(g19943,g7562,g18976);
  and AND2_1996(g19944,g3028,g18258);
  and AND2_1997(g19949,g5293,g18278);
  and AND2_1998(g19952,g2760,g18987);
  and AND2_1999(g19953,g7566,g18334);
  and AND3_90(II26416,g18553,g18491,g18431);
  and AND3_91(g19970,g18354,g18276,II26416);
  and AND2_2000(g19971,g5327,g18355);
  and AND2_2001(g19976,g5330,g18371);
  and AND3_92(II26432,g18277,g18189,g18090);
  and AND3_93(g19982,g17992,g17913,II26432);
  and AND2_2002(g19983,g5352,g18432);
  and AND3_94(II26440,g18603,g18555,g18504);
  and AND3_95(g20000,g18449,g18369,II26440);
  and AND2_2003(g20001,g5355,g18450);
  and AND2_2004(g20006,g5358,g18466);
  and AND2_2005(g20011,g18063,g3113);
  and AND2_2006(g20012,g16804,g3135);
  and AND2_2007(g20013,g17720,g12848);
  and AND2_2008(g20014,g7615,g16749);
  and AND3_96(II26464,g18370,g18296,g18206);
  and AND3_97(g20020,g18109,g18024,II26464);
  and AND2_2009(g20021,g5369,g18505);
  and AND3_98(II26472,g18635,g18605,g18568);
  and AND3_99(g20038,g18522,g18464,II26472);
  and AND2_2010(g20039,g5372,g18523);
  and AND2_2011(g20044,g5375,g18539);
  and AND2_2012(g20048,g16749,g3127);
  and AND2_2013(g20049,g17878,g3155);
  and AND2_2014(g20050,g18070,g3161);
  and AND2_2015(g20051,g18063,g3114);
  and AND2_2016(g20052,g16804,g3134);
  and AND2_2017(g20053,g17720,g12875);
  and AND3_100(II26500,g18465,g18389,g18313);
  and AND3_101(g20062,g18225,g18141,II26500);
  and AND2_2018(g20063,g5382,g18569);
  and AND3_102(II26508,g18644,g18637,g18618);
  and AND3_103(g20080,g18586,g18537,II26508);
  and AND2_2019(g20081,g5385,g18587);
  and AND2_2020(g20084,g17969,g3158);
  and AND2_2021(g20085,g18170,g3164);
  and AND2_2022(g20086,g18337,g3170);
  and AND2_2023(g20087,g16749,g7574);
  and AND2_2024(g20088,g16836,g3147);
  and AND2_2025(g20089,g17969,g9160);
  and AND2_2026(g20090,g18063,g3120);
  and AND2_2027(g20091,g16804,g3136);
  and AND2_2028(g20092,g16749,g7603);
  and AND3_104(II26525,g18656,g18670,g18692);
  and AND4_61(g20093,g13657,g13677,g13750,II26525);
  and AND3_105(II26528,g18656,g14837,g13657);
  and AND3_106(g20094,g13677,g13706,II26528);
  and AND3_107(II26541,g18538,g18484,g18406);
  and AND3_108(g20103,g18332,g18257,II26541);
  and AND2_2029(g20104,g5391,g18619);
  and AND2_2030(g20106,g18261,g3167);
  and AND2_2031(g20107,g18415,g3173);
  and AND2_2032(g20108,g18543,g3179);
  and AND2_2033(g20109,g17878,g9504);
  and AND2_2034(g20110,g18070,g9286);
  and AND2_2035(g20111,g18261,g9884);
  and AND2_2036(g20112,g16749,g3132);
  and AND2_2037(g20113,g16836,g3142);
  and AND2_2038(g20114,g17969,g9755);
  and AND2_2039(g20115,g16804,g3139);
  and AND3_109(II26558,g14776,g18670,g18720);
  and AND4_62(g20116,g16142,g13677,g13706,II26558);
  and AND3_110(II26561,g14776,g18720,g13657);
  and AND3_111(g20117,g16189,g13706,II26561);
  and AND3_112(II26564,g18679,g18699,g18728);
  and AND4_63(g20118,g13687,g13714,g13791,II26564);
  and AND3_113(II26567,g18679,g14910,g13687);
  and AND3_114(g20119,g13714,g13756,II26567);
  and AND2_2040(g20131,g18486,g3176);
  and AND2_2041(g20132,g18593,g3182);
  and AND2_2042(g20133,g18170,g9505);
  and AND2_2043(g20134,g18337,g9506);
  and AND2_2044(g20135,g18486,g9885);
  and AND2_2045(g20136,g17878,g9423);
  and AND2_2046(g20137,g18070,g9226);
  and AND2_2047(g20138,g18261,g9756);
  and AND2_2048(g20139,g16836,g3151);
  and AND3_115(g20144,g16679,g16884,g16665);
  and AND4_64(g20145,g14776,g18670,g16142,g16189);
  and AND3_116(II26590,g14811,g18699,g18758);
  and AND4_65(g20146,g16201,g13714,g13756,II26590);
  and AND3_117(II26593,g14811,g18758,g13687);
  and AND3_118(g20147,g16254,g13756,II26593);
  and AND3_119(II26596,g18708,g18735,g18765);
  and AND4_66(g20148,g13724,g13764,g13819,II26596);
  and AND3_120(II26599,g18708,g14991,g13724);
  and AND3_121(g20149,g13764,g13797,II26599);
  and AND2_2049(g20156,g16809,g3185);
  and AND2_2050(g20157,g18415,g9287);
  and AND2_2051(g20158,g18543,g9886);
  and AND2_2052(g20159,g16809,g9288);
  and AND2_2053(g20160,g18170,g9424);
  and AND2_2054(g20161,g18337,g9426);
  and AND2_2055(g20162,g18486,g9757);
  and AND3_122(II26615,g14797,g18692,g13657);
  and AND3_123(g20177,g13677,g13750,II26615);
  and AND3_124(g20182,g16705,g16913,g16686);
  and AND4_67(g20183,g14811,g18699,g16201,g16254);
  and AND3_125(II26621,g14863,g18735,g18789);
  and AND4_68(g20184,g16266,g13764,g13797,II26621);
  and AND3_126(II26624,g14863,g18789,g13724);
  and AND3_127(g20185,g16313,g13797,II26624);
  and AND3_128(II26627,g18744,g18772,g18796);
  and AND4_69(g20186,g13774,g13805,g13840,II26627);
  and AND3_129(II26630,g18744,g15080,g13774);
  and AND3_130(g20187,g13805,g13825,II26630);
  and AND2_2056(g20188,g18593,g9425);
  and AND2_2057(g20189,g16825,g9289);
  and AND2_2058(g20190,g18415,g9227);
  and AND2_2059(g20191,g18543,g9758);
  and AND2_2060(g20192,g16809,g9228);
  and AND3_131(II26639,g18656,g18670,g16142);
  and AND3_132(g20197,g13677,g13706,II26639);
  and AND3_133(II26645,g14849,g18728,g13687);
  and AND3_134(g20211,g13714,g13791,II26645);
  and AND3_135(g20216,g16736,g16943,g16712);
  and AND4_70(g20217,g14863,g18735,g16266,g16313);
  and AND3_136(II26651,g14936,g18772,g18815);
  and AND4_71(g20218,g16325,g13805,g13825,II26651);
  and AND3_137(II26654,g14936,g18815,g13774);
  and AND3_138(g20219,g16371,g13825,II26654);
  and AND2_2061(g20220,g18593,g9355);
  and AND2_2062(g20221,g16825,g10099);
  and AND4_72(g20222,g18656,g18720,g13657,g16293);
  and AND3_139(II26661,g18679,g18699,g16201);
  and AND3_140(g20227,g13714,g13756,II26661);
  and AND3_141(II26667,g14922,g18765,g13724);
  and AND3_142(g20241,g13764,g13819,II26667);
  and AND3_143(g20246,g16778,g16974,g16743);
  and AND4_73(g20247,g14936,g18772,g16325,g16371);
  and AND3_144(g20248,g18656,g14837,g16293);
  and AND4_74(g20249,g18679,g18758,g13687,g16351);
  and AND3_145(II26676,g18708,g18735,g16266);
  and AND3_146(g20254,g13764,g13797,II26676);
  and AND3_147(II26682,g15003,g18796,g13774);
  and AND3_148(g20268,g13805,g13840,II26682);
  and AND4_75(g20270,g14797,g18692,g13657,g16243);
  and AND3_149(g20271,g18679,g14910,g16351);
  and AND4_76(g20272,g18708,g18789,g13724,g16395);
  and AND3_150(II26690,g18744,g18772,g16325);
  and AND3_151(g20277,g13805,g13825,II26690);
  and AND3_152(II26695,g18670,g18692,g16142);
  and AND3_153(g20280,g13677,g16243,II26695);
  and AND4_77(g20282,g14849,g18728,g13687,g16302);
  and AND3_154(g20283,g18708,g14991,g16395);
  and AND4_78(g20284,g18744,g18815,g13774,g16433);
  and AND2_2063(g20285,g16846,g8103);
  and AND3_155(II26708,g18699,g18728,g16201);
  and AND3_156(g20291,g13714,g16302,II26708);
  and AND4_79(g20293,g14922,g18765,g13724,g16360);
  and AND3_157(g20294,g18744,g15080,g16433);
  and AND3_158(II26726,g18735,g18765,g16266);
  and AND3_159(g20307,g13764,g16360,II26726);
  and AND4_80(g20309,g15003,g18796,g13774,g16404);
  and AND3_160(II26745,g18772,g18796,g16325);
  and AND3_161(g20326,g13805,g16404,II26745);
  and AND2_2064(g20460,g17351,g13644);
  and AND2_2065(g20472,g17314,g13669);
  and AND2_2066(g20480,g17313,g11827);
  and AND2_2067(g20486,g17281,g11859);
  and AND2_2068(g20492,g17258,g11894);
  and AND2_2069(g20499,g17648,g11933);
  and AND2_2070(g20502,g17566,g11973);
  and AND2_2071(g20503,g17507,g13817);
  and AND2_2072(g20506,g17499,g12025);
  and AND2_2073(g20512,g17445,g13836);
  and AND2_2074(g20525,g17394,g13849);
  and AND4_81(g20538,g18656,g14837,g13657,g16189);
  and AND2_2075(g20640,g4809,g19064);
  and AND2_2076(g20647,g5888,g19075);
  and AND2_2077(g20665,g4985,g19081);
  and AND2_2078(g20809,g5712,g19113);
  and AND2_2079(g20826,g5770,g19118);
  and AND2_2080(g20836,g5829,g19125);
  and AND2_2081(g20840,g5885,g19132);
  and AND3_162(g21049,g20016,g14079,g14165);
  and AND2_2082(g21067,g20193,g12030);
  and AND3_163(g21068,g20058,g14194,g14280);
  and AND2_2083(g21077,g20223,g12094);
  and AND3_164(g21078,g20099,g14309,g14402);
  and AND3_165(g21085,g19484,g14158,g19001);
  and AND2_2084(g21086,g20193,g12142);
  and AND2_2085(g21091,g20250,g12166);
  and AND3_166(g21092,g20124,g14431,g14514);
  and AND3_167(g21097,g19505,g14273,g16507);
  and AND2_2086(g21098,g20223,g12204);
  and AND2_2087(g21103,g20273,g12228);
  and AND3_168(g21107,g19444,g17893,g14079);
  and AND3_169(g21111,g19524,g14395,g16529);
  and AND2_2088(g21112,g20250,g12259);
  and AND2_2089(g21121,g20054,g14244);
  and AND2_2090(g21122,g20140,g12279);
  and AND2_2091(g21123,g19970,g19982);
  and AND3_170(g21124,g19471,g18004,g14194);
  and AND3_171(g21128,g19534,g14507,g16560);
  and AND2_2092(g21129,g20273,g12302);
  and AND3_172(II27695,g19318,g19300,g19286);
  and AND3_173(g21136,g19271,g19261,II27695);
  and AND2_2093(g21137,g5750,g19272);
  and AND2_2094(g21138,g19484,g14347);
  and AND2_2095(g21140,g20095,g14366);
  and AND2_2096(g21141,g20178,g12315);
  and AND2_2097(g21142,g20000,g20020);
  and AND3_174(g21143,g19494,g18121,g14309);
  and AND3_175(II27711,g19262,g19414,g19386);
  and AND3_176(g21152,g19357,g19334,II27711);
  and AND3_177(g21153,g20054,g16543,g16501);
  and AND2_2098(g21154,g20193,g12333);
  and AND2_2099(g21155,g20140,g12336);
  and AND3_178(II27717,g19345,g19321,g19304);
  and AND3_179(g21156,g19290,g19276,II27717);
  and AND2_2100(g21157,g5809,g19291);
  and AND2_2101(g21158,g19505,g14459);
  and AND2_2102(g21160,g20120,g14478);
  and AND2_2103(g21161,g20212,g12343);
  and AND2_2104(g21162,g20038,g20062);
  and AND3_180(g21163,g19515,g18237,g14431);
  and AND3_181(II27733,g19277,g19451,g19416);
  and AND3_182(g21172,g19389,g19368,II27733);
  and AND3_183(g21173,g20095,g16575,g16523);
  and AND2_2105(g21174,g20223,g12363);
  and AND2_2106(g21175,g20178,g12366);
  and AND3_184(II27739,g19379,g19348,g19325);
  and AND3_185(g21176,g19308,g19295,II27739);
  and AND2_2107(g21177,g5865,g19309);
  and AND2_2108(g21178,g19524,g14546);
  and AND2_2109(g21180,g20150,g14565);
  and AND2_2110(g21181,g20242,g12373);
  and AND2_2111(g21182,g20080,g20103);
  and AND2_2112(g21188,g20140,g12379);
  and AND3_186(II27755,g19296,g19478,g19453);
  and AND3_187(g21192,g19419,g19400,II27755);
  and AND3_188(g21193,g20120,g16599,g16554);
  and AND2_2113(g21194,g20250,g12382);
  and AND2_2114(g21195,g20212,g12385);
  and AND3_189(II27761,g19411,g19382,g19352);
  and AND3_190(g21196,g19329,g19313,II27761);
  and AND2_2115(g21197,g5912,g19330);
  and AND2_2116(g21198,g19534,g14601);
  and AND2_2117(g21203,g20178,g12409);
  and AND3_191(II27772,g19314,g19501,g19480);
  and AND3_192(g21207,g19456,g19430,II27772);
  and AND3_193(g21208,g20150,g16619,g16586);
  and AND2_2118(g21209,g20273,g12412);
  and AND2_2119(g21210,g20242,g12415);
  and AND2_2120(g21218,g20212,g12421);
  and AND2_2121(g21226,g20242,g12426);
  and AND3_194(g21229,g19578,g14797,g16665);
  and AND3_195(g21234,g19608,g14849,g16686);
  and AND3_196(g21243,g19641,g14922,g16712);
  and AND2_2122(g21245,g20299,g14837);
  and AND3_197(g21251,g19681,g15003,g16743);
  and AND2_2123(g21252,g19578,g14895);
  and AND2_2124(g21254,g20318,g14910);
  and AND3_198(g21259,g20299,g16722,g16682);
  and AND2_2125(g21260,g19608,g14976);
  and AND2_2126(g21262,g20337,g14991);
  and AND3_199(g21267,g20318,g16764,g16708);
  and AND2_2127(g21268,g19641,g15065);
  and AND2_2128(g21270,g20357,g15080);
  and AND3_200(g21276,g20337,g16791,g16739);
  and AND2_2129(g21277,g19681,g15161);
  and AND3_201(g21283,g20357,g16820,g16781);
  and AND2_2130(g21284,g9356,g20269);
  and AND2_2131(g21290,g9356,g20278);
  and AND2_2132(g21291,g9293,g20279);
  and AND2_2133(g21292,g9453,g20281);
  and AND2_2134(g21298,g9356,g20286);
  and AND2_2135(g21299,g9293,g20287);
  and AND2_2136(g21300,g9232,g20288);
  and AND2_2137(g21301,g9453,g20289);
  and AND2_2138(g21302,g9374,g20290);
  and AND2_2139(g21303,g9595,g20292);
  and AND2_2140(g21304,g9293,g20296);
  and AND2_2141(g21305,g9232,g20297);
  and AND2_2142(g21306,g9187,g20298);
  and AND2_2143(g21307,g9453,g20302);
  and AND2_2144(g21308,g9374,g20303);
  and AND2_2145(g21309,g9310,g20304);
  and AND2_2146(g21310,g9595,g20305);
  and AND2_2147(g21311,g9471,g20306);
  and AND2_2148(g21312,g9737,g20308);
  and AND2_2149(g21313,g9232,g20311);
  and AND2_2150(g21314,g9187,g20312);
  and AND2_2151(g21315,g9161,g20313);
  and AND2_2152(g21319,g9374,g20315);
  and AND2_2153(g21320,g9310,g20316);
  and AND2_2154(g21321,g9248,g20317);
  and AND2_2155(g21322,g9595,g20321);
  and AND2_2156(g21323,g9471,g20322);
  and AND2_2157(g21324,g9391,g20323);
  and AND2_2158(g21325,g9737,g20324);
  and AND2_2159(g21326,g9613,g20325);
  and AND2_2160(g21328,g9187,g20327);
  and AND2_2161(g21329,g9161,g20328);
  and AND2_2162(g21330,g9150,g20329);
  and AND2_2163(g21334,g9310,g20330);
  and AND2_2164(g21335,g9248,g20331);
  and AND2_2165(g21336,g9203,g20332);
  and AND2_2166(g21337,g9471,g20334);
  and AND2_2167(g21338,g9391,g20335);
  and AND2_2168(g21339,g9326,g20336);
  and AND2_2169(g21340,g9737,g20340);
  and AND2_2170(g21341,g9613,g20341);
  and AND2_2171(g21342,g9488,g20342);
  and AND2_2172(g21343,g9161,g20344);
  and AND2_2173(g21344,g9150,g20345);
  and AND2_2174(g21345,g15096,g20346);
  and AND2_2175(g21349,g9248,g20347);
  and AND2_2176(g21350,g9203,g20348);
  and AND2_2177(g21351,g9174,g20349);
  and AND2_2178(g21352,g9391,g20350);
  and AND2_2179(g21353,g9326,g20351);
  and AND2_2180(g21354,g9264,g20352);
  and AND2_2181(g21355,g9613,g20354);
  and AND2_2182(g21356,g9488,g20355);
  and AND2_2183(g21357,g9407,g20356);
  and AND2_2184(g21360,g9507,g20361);
  and AND2_2185(g21361,g9150,g20362);
  and AND2_2186(g21362,g15096,g20363);
  and AND2_2187(g21363,g15022,g20364);
  and AND2_2188(g21367,g9203,g20366);
  and AND2_2189(g21368,g9174,g20367);
  and AND2_2190(g21369,g15188,g20368);
  and AND2_2191(g21370,g9326,g20369);
  and AND2_2192(g21371,g9264,g20370);
  and AND2_2193(g21372,g9216,g20371);
  and AND2_2194(g21373,g9488,g20372);
  and AND2_2195(g21374,g9407,g20373);
  and AND2_2196(g21375,g9342,g20374);
  and AND2_2197(g21378,g9507,g20378);
  and AND2_2198(g21379,g9427,g20379);
  and AND2_2199(g21380,g15096,g20380);
  and AND2_2200(g21381,g15022,g20381);
  and AND2_2201(g21388,g6201,g19657);
  and AND2_2202(g21389,g9649,g20384);
  and AND2_2203(g21390,g9174,g20385);
  and AND2_2204(g21391,g15188,g20386);
  and AND2_2205(g21392,g15118,g20387);
  and AND2_2206(g21393,g9264,g20389);
  and AND2_2207(g21394,g9216,g20390);
  and AND2_2208(g21395,g15274,g20391);
  and AND2_2209(g21396,g9407,g20392);
  and AND2_2210(g21397,g9342,g20393);
  and AND2_2211(g21398,g9277,g20394);
  and AND2_2212(g21401,g9507,g20397);
  and AND2_2213(g21402,g9427,g20398);
  and AND2_2214(g21403,g15022,g20399);
  and AND2_2215(g21410,g6363,g20402);
  and AND2_2216(g21411,g9649,g20403);
  and AND2_2217(g21412,g9569,g20404);
  and AND2_2218(g21413,g15188,g20405);
  and AND2_2219(g21414,g15118,g20406);
  and AND2_2220(g21418,g6290,g19705);
  and AND2_2221(g21419,g9795,g20409);
  and AND2_2222(g21420,g9216,g20410);
  and AND2_2223(g21421,g15274,g20411);
  and AND2_2224(g21422,g15210,g20412);
  and AND2_2225(g21423,g9342,g20414);
  and AND2_2226(g21424,g9277,g20415);
  and AND2_2227(g21425,g15366,g20416);
  and AND2_2228(g21428,g9427,g20420);
  and AND2_2229(g21438,g9649,g20422);
  and AND2_2230(g21439,g9569,g20423);
  and AND2_2231(g21440,g15118,g20424);
  and AND2_2232(g21444,g6568,g20427);
  and AND2_2233(g21445,g9795,g20428);
  and AND2_2234(g21446,g9711,g20429);
  and AND2_2235(g21447,g15274,g20430);
  and AND2_2236(g21448,g15210,g20431);
  and AND2_2237(g21452,g6427,g19749);
  and AND2_2238(g21453,g9941,g20434);
  and AND2_2239(g21454,g9277,g20435);
  and AND2_2240(g21455,g15366,g20436);
  and AND2_2241(g21456,g15296,g20437);
  and AND2_2242(g21476,g9569,g20442);
  and AND2_2243(g21480,g9795,g20444);
  and AND2_2244(g21481,g9711,g20445);
  and AND2_2245(g21482,g15210,g20446);
  and AND2_2246(g21486,g6832,g20449);
  and AND2_2247(g21487,g9941,g20450);
  and AND2_2248(g21488,g9857,g20451);
  and AND2_2249(g21489,g15366,g20452);
  and AND2_2250(g21490,g15296,g20453);
  and AND2_2251(g21494,g6632,g19792);
  and AND2_2252(g21497,g3006,g20456);
  and AND2_2253(g21517,g9711,g20461);
  and AND2_2254(g21521,g9941,g20463);
  and AND2_2255(g21522,g9857,g20464);
  and AND2_2256(g21523,g15296,g20465);
  and AND2_2257(g21527,g7134,g20468);
  and AND3_202(II28068,g17802,g18265,g17882);
  and AND4_82(g21533,g17724,g18179,g19799,II28068);
  and AND2_2258(g21553,g9857,g20476);
  and AND3_203(II28096,g13907,g14238,g13946);
  and AND4_83(g21564,g13886,g14153,g19799,II28096);
  and AND3_204(II28103,g17914,g18358,g17993);
  and AND4_84(g21569,g17825,g18286,g19843,II28103);
  and AND2_2259(g21589,g3002,g19890);
  and AND3_205(g21593,g16498,g19484,g14071);
  and AND3_206(II28126,g13963,g14360,g14016);
  and AND4_85(g21597,g13927,g14268,g19843,II28126);
  and AND3_207(II28133,g18025,g18453,g18110);
  and AND4_86(g21602,g17937,g18379,g19876,II28133);
  and AND2_2260(g21610,g7522,g20490);
  and AND2_2261(g21611,g7471,g19915);
  and AND3_208(g21622,g16520,g19505,g14186);
  and AND3_209(II28155,g14033,g14472,g14107);
  and AND4_87(g21626,g13983,g14390,g19876,II28155);
  and AND3_210(II28162,g18142,g18526,g18226);
  and AND4_88(g21631,g18048,g18474,g19907,II28162);
  and AND2_2262(g21635,g7549,g20496);
  and AND2_2263(g21639,g3398,g20500);
  and AND3_211(g21650,g16551,g19524,g14301);
  and AND3_212(II28181,g14124,g14559,g14222);
  and AND4_89(g21654,g14053,g14502,g19907,II28181);
  and AND2_2264(g21658,g2896,g20501);
  and AND2_2265(g21666,g3398,g20504);
  and AND2_2266(g21670,g3554,g20505);
  and AND3_213(g21681,g16583,g19534,g14423);
  and AND2_2267(g21687,g3398,g20516);
  and AND2_2268(g21695,g3554,g20517);
  and AND2_2269(g21699,g3710,g20518);
  and AND2_2270(g21707,g2892,g19978);
  and AND2_2271(g21723,g3554,g20534);
  and AND2_2272(g21731,g3710,g20535);
  and AND2_2273(g21735,g3866,g20536);
  and AND2_2274(g21749,g3710,g20553);
  and AND2_2275(g21757,g3866,g20554);
  and AND2_2276(g21758,g7607,g20045);
  and AND2_2277(g21773,g3866,g19078);
  and AND3_214(g21805,g16679,g19578,g14776);
  and AND3_215(g21812,g16705,g19608,g14811);
  and AND3_216(g21818,g16736,g19641,g14863);
  and AND3_217(g21822,g16778,g19681,g14936);
  and AND2_2278(g21891,g19302,g11749);
  and AND2_2279(g21892,g19288,g13011);
  and AND2_2280(g21899,g19323,g11749);
  and AND2_2281(g21900,g19306,g13011);
  and AND2_2282(g21906,g5715,g20513);
  and AND2_2283(g21911,g19350,g11749);
  and AND2_2284(g21912,g19327,g13011);
  and AND2_2285(g21913,g4456,g20519);
  and AND2_2286(g21920,g5773,g20531);
  and AND2_2287(g21925,g19384,g11749);
  and AND2_2288(g21926,g19354,g13011);
  and AND2_2289(g21931,g4632,g20539);
  and AND2_2290(g21938,g5832,g20550);
  and AND2_2291(g21990,g291,g21187);
  and AND2_2292(g22004,g978,g21202);
  and AND2_2293(g22015,g1672,g21217);
  and AND2_2294(g22020,g2366,g21225);
  and AND3_218(II28582,g19141,g21133,g21116);
  and AND4_90(g22036,g21104,g21095,g21084,II28582);
  and AND3_219(II28594,g21167,g21147,g21134);
  and AND4_91(g22046,g21117,g21105,g21096,II28594);
  and AND3_220(II28609,g21183,g21168,g21148);
  and AND4_92(g22062,g21135,g21118,g21106,II28609);
  and AND2_2295(g22187,g21564,g20986);
  and AND2_2296(g22196,g21597,g21012);
  and AND2_2297(g22201,g21271,g16881);
  and AND2_2298(g22202,g21626,g21036);
  and AND2_2299(g22206,g21895,g11976);
  and AND2_2300(g22207,g21278,g16910);
  and AND2_2301(g22208,g21654,g21057);
  and AND2_2302(g22211,g21661,g12027);
  and AND2_2303(g22214,g21907,g12045);
  and AND2_2304(g22215,g21285,g16940);
  and AND2_2305(g22220,g21690,g12091);
  and AND2_2306(g22223,g21921,g12109);
  and AND2_2307(g22224,g21293,g16971);
  and AND2_2308(g22228,g21716,g12136);
  and AND2_2309(g22229,g21661,g12139);
  and AND2_2310(g22235,g21726,g12163);
  and AND2_2311(g22238,g21939,g12181);
  and AND2_2312(g22244,g21742,g12198);
  and AND2_2313(g22245,g21690,g12201);
  and AND2_2314(g22250,g21752,g12225);
  and AND2_2315(g22254,g21716,g12239);
  and AND2_2316(g22255,g21661,g12242);
  and AND2_2317(g22264,g21766,g12253);
  and AND2_2318(g22265,g21726,g12256);
  and AND2_2319(g22270,g92,g21529);
  and AND2_2320(g22272,g21742,g12282);
  and AND2_2321(g22273,g21690,g12285);
  and AND2_2322(g22281,g21782,g12296);
  and AND2_2323(g22282,g21752,g12299);
  and AND2_2324(g22285,g21716,g12312);
  and AND2_2325(g22289,g780,g21565);
  and AND2_2326(g22291,g21766,g12318);
  and AND2_2327(g22292,g21726,g12321);
  and AND2_2328(g22305,g21742,g12340);
  and AND2_2329(g22309,g1466,g21598);
  and AND2_2330(g22311,g21782,g12346);
  and AND2_2331(g22312,g21752,g12349);
  and AND2_2332(g22333,g21766,g12370);
  and AND2_2333(g22337,g2160,g21627);
  and AND2_2334(g22340,g88,g21184);
  and AND2_2335(g22358,g21782,g12389);
  and AND2_2336(g22363,g776,g21199);
  and AND2_2337(g22383,g1462,g21214);
  and AND2_2338(g22398,g2156,g21222);
  and AND2_2339(g22483,g646,g21861);
  and AND2_2340(g22515,g13873,g21382);
  and AND2_2341(g22516,g20885,g17442);
  and AND2_2342(g22517,g21895,g12608);
  and AND2_2343(g22526,g1332,g21867);
  and AND2_2344(g22546,g13886,g21404);
  and AND2_2345(g22555,g13895,g21415);
  and AND2_2346(g22556,g20904,g17523);
  and AND2_2347(g22557,g21907,g12654);
  and AND2_2348(g22566,g2026,g21872);
  and AND2_2349(g22577,g13907,g21429);
  and AND2_2350(g22581,g21895,g12699);
  and AND2_2351(g22587,g13927,g21441);
  and AND2_2352(g22595,g13936,g21449);
  and AND2_2353(g22596,g20928,g17613);
  and AND2_2354(g22597,g21921,g12708);
  and AND2_2355(g22606,g2720,g21876);
  and AND2_2356(g22607,g13946,g21458);
  and AND2_2357(g22610,g660,g21473);
  and AND2_2358(g22614,g13963,g21477);
  and AND2_2359(g22618,g21907,g12756);
  and AND2_2360(g22624,g13983,g21483);
  and AND2_2361(g22632,g13992,g21491);
  and AND2_2362(g22633,g20956,g17710);
  and AND2_2363(g22634,g21939,g12765);
  and AND2_2364(g22637,g20841,g10927);
  and AND2_2365(g22638,g14001,g21498);
  and AND2_2366(g22643,g14016,g21505);
  and AND2_2367(g22646,g1346,g21514);
  and AND2_2368(g22650,g14033,g21518);
  and AND2_2369(g22654,g21921,g12798);
  and AND2_2370(g22660,g14053,g21524);
  and AND2_2371(g22665,g20920,g6153);
  and AND2_2372(g22666,g21825,g20014);
  and AND2_2373(g22667,g14062,g21530);
  and AND2_2374(g22674,g14092,g21537);
  and AND2_2375(g22679,g14107,g21541);
  and AND2_2376(g22682,g2040,g21550);
  and AND2_2377(g22686,g14124,g21554);
  and AND2_2378(g22690,g21939,g12837);
  and AND2_2379(g22699,g7338,g21883);
  and AND2_2380(g22700,g7146,g21558);
  and AND2_2381(g22701,g18174,g21561);
  and AND2_2382(g22707,g14177,g21566);
  and AND2_2383(g22714,g14207,g21573);
  and AND2_2384(g22719,g14222,g21577);
  and AND2_2385(g22722,g2734,g21586);
  and AND2_2386(g22726,g3036,g21886);
  and AND2_2387(g22727,g14238,g21590);
  and AND2_2388(g22732,g18281,g21594);
  and AND2_2389(g22738,g14292,g21599);
  and AND2_2390(g22745,g14322,g21606);
  and AND2_2391(g22754,g14342,g21612);
  and AND2_2392(g22759,g14360,g21619);
  and AND2_2393(g22764,g18374,g21623);
  and AND2_2394(g22770,g14414,g21628);
  and AND2_2395(g22788,g14454,g21640);
  and AND2_2396(g22793,g14472,g21647);
  and AND2_2397(g22798,g18469,g21651);
  and AND2_2398(g22804,g2920,g21655);
  and AND2_2399(g22830,g14541,g21671);
  and AND2_2400(g22835,g14559,g21678);
  and AND2_2401(g22841,g7583,g21902);
  and AND2_2402(g22842,g3032,g21682);
  and AND2_2403(g22869,g14596,g21700);
  and AND2_2404(g22874,g7587,g21708);
  and AND2_2405(g22906,g2924,g21927);
  and AND2_2406(g22984,g16840,g21400);
  and AND2_2407(g23104,g20842,g15859);
  and AND2_2408(g23106,g5857,g21050);
  and AND2_2409(g23118,g20850,g15890);
  and AND2_2410(g23119,g5904,g21069);
  and AND2_2411(g23127,g20858,g15923);
  and AND2_2412(g23128,g5943,g21079);
  and AND2_2413(g23138,g20866,g15952);
  and AND2_2414(g23139,g5977,g21093);
  and AND2_2415(g23409,g21533,g22408);
  and AND2_2416(g23414,g21569,g22421);
  and AND2_2417(g23419,g22755,g19577);
  and AND2_2418(g23423,g21602,g22443);
  and AND2_2419(g23428,g22789,g19607);
  and AND2_2420(g23432,g21631,g22476);
  and AND2_2421(g23434,g22831,g19640);
  and AND2_2422(g23440,g22870,g19680);
  and AND2_2423(g23451,g18552,g22547);
  and AND2_2424(g23458,g18602,g22588);
  and AND2_2425(g23462,g17988,g22609);
  and AND2_2426(g23467,g18634,g22625);
  and AND2_2427(g23471,g18105,g22645);
  and AND2_2428(g23476,g18643,g22661);
  and AND2_2429(g23483,g22945,g8847);
  and AND2_2430(g23484,g18221,g22681);
  and AND2_2431(g23494,g18328,g22721);
  and AND2_2432(g23496,g5802,g22300);
  and AND2_2433(g23510,g5890,g22753);
  and AND2_2434(g23512,g5858,g22328);
  and AND2_2435(g23525,g5929,g22787);
  and AND2_2436(g23527,g5905,g22353);
  and AND2_2437(g23536,g5963,g22829);
  and AND2_2438(g23538,g5944,g22376);
  and AND2_2439(g23544,g5992,g22868);
  and AND2_2440(g23547,g8062,g22405);
  and AND2_2441(g23550,g8132,g22409);
  and AND2_2442(g23551,g8135,g22412);
  and AND2_2443(g23552,g6136,g22415);
  and AND2_2444(g23554,g8147,g22418);
  and AND2_2445(g23558,g8200,g22422);
  and AND2_2446(g23559,g8203,g22425);
  and AND2_2447(g23560,g8206,g22428);
  and AND2_2448(g23563,g8218,g22431);
  and AND2_2449(g23564,g8221,g22434);
  and AND2_2450(g23565,g6146,g22437);
  and AND2_2451(g23567,g8233,g22440);
  and AND2_2452(g23571,g3931,g22445);
  and AND2_2453(g23572,g3934,g22448);
  and AND2_2454(g23573,g3937,g22451);
  and AND2_2455(g23577,g3957,g22455);
  and AND2_2456(g23578,g3960,g22458);
  and AND2_2457(g23579,g3963,g22461);
  and AND2_2458(g23582,g3975,g22464);
  and AND2_2459(g23583,g3978,g22467);
  and AND2_2460(g23584,g6167,g22470);
  and AND2_2461(g23586,g3990,g22473);
  and AND2_2462(g23590,g4009,g22477);
  and AND2_2463(g23591,g4012,g22480);
  and AND2_2464(g23592,g17640,g22986);
  and AND2_2465(g23593,g22845,g20365);
  and AND2_2466(g23598,g4038,g22484);
  and AND2_2467(g23599,g4041,g22487);
  and AND2_2468(g23600,g4044,g22490);
  and AND2_2469(g23604,g4064,g22494);
  and AND2_2470(g23605,g4067,g22497);
  and AND2_2471(g23606,g4070,g22500);
  and AND2_2472(g23609,g4082,g22503);
  and AND2_2473(g23610,g4085,g22506);
  and AND2_2474(g23611,g6194,g22509);
  and AND2_2475(g23615,g4107,g22512);
  and AND2_2476(g23616,g17724,g22988);
  and AND2_2477(g23617,g22810,g20382);
  and AND2_2478(g23618,g22608,g20383);
  and AND2_2479(g23622,g4136,g22520);
  and AND2_2480(g23623,g4139,g22523);
  and AND2_2481(g23624,g17741,g22989);
  and AND2_2482(g23625,g22880,g20388);
  and AND2_2483(g23630,g4165,g22527);
  and AND2_2484(g23631,g4168,g22530);
  and AND2_2485(g23632,g4171,g22533);
  and AND2_2486(g23636,g4191,g22537);
  and AND2_2487(g23637,g4194,g22540);
  and AND2_2488(g23638,g4197,g22543);
  and AND2_2489(g23639,g21825,g22805);
  and AND2_2490(g23643,g17802,g22991);
  and AND2_2491(g23659,g22784,g17500);
  and AND2_2492(g23664,g4246,g22552);
  and AND2_2493(g23665,g17825,g22995);
  and AND2_2494(g23666,g22851,g20407);
  and AND2_2495(g23667,g22644,g20408);
  and AND2_2496(g23671,g4275,g22560);
  and AND2_2497(g23672,g4278,g22563);
  and AND2_2498(g23673,g17842,g22996);
  and AND2_2499(g23674,g22915,g20413);
  and AND2_2500(g23679,g4304,g22567);
  and AND2_2501(g23680,g4307,g22570);
  and AND2_2502(g23681,g4310,g22573);
  and AND2_2503(g23686,g17882,g22998);
  and AND2_2504(g23687,g22668,g17570);
  and AND2_2505(g23689,g6513,g23001);
  and AND2_2506(g23693,g17914,g23002);
  and AND2_2507(g23709,g22826,g17591);
  and AND2_2508(g23714,g4401,g22592);
  and AND2_2509(g23715,g17937,g23006);
  and AND2_2510(g23716,g22886,g20432);
  and AND2_2511(g23717,g22680,g20433);
  and AND2_2512(g23721,g4430,g22600);
  and AND2_2513(g23722,g4433,g22603);
  and AND2_2514(g23723,g17954,g23007);
  and AND2_2515(g23724,g22940,g20438);
  and AND2_2516(g23726,g21825,g22843);
  and AND2_2517(g23734,g17974,g23008);
  and AND2_2518(g23735,g22949,g9450);
  and AND2_2519(g23740,g17993,g23012);
  and AND2_2520(g23741,g22708,g17667);
  and AND2_2521(g23743,g6777,g23015);
  and AND2_2522(g23747,g18025,g23016);
  and AND2_2523(g23763,g22865,g17688);
  and AND2_2524(g23768,g4570,g22629);
  and AND2_2525(g23769,g18048,g23020);
  and AND2_2526(g23770,g22921,g20454);
  and AND2_2527(g23771,g22720,g20455);
  and AND2_2528(g23772,g21825,g22875);
  and AND2_2529(g23776,g18074,g23021);
  and AND2_2530(g23777,g22949,g9528);
  and AND2_2531(g23778,g22954,g9531);
  and AND2_2532(g23789,g18091,g23024);
  and AND2_2533(g23790,g22958,g9592);
  and AND2_2534(g23795,g18110,g23028);
  and AND2_2535(g23796,g22739,g17767);
  and AND2_2536(g23798,g7079,g23031);
  and AND2_2537(g23802,g18142,g23032);
  and AND2_2538(g23818,g22900,g17788);
  and AND2_2539(g23820,g3013,g23036);
  and AND2_2540(g23822,g14148,g23037);
  and AND2_2541(g23824,g22949,g9641);
  and AND2_2542(g23825,g22954,g9644);
  and AND2_2543(g23829,g18190,g23038);
  and AND2_2544(g23830,g22958,g9670);
  and AND2_2545(g23831,g22962,g9673);
  and AND2_2546(g23842,g18207,g23041);
  and AND2_2547(g23843,g22966,g9734);
  and AND2_2548(g23848,g18226,g23045);
  and AND2_2549(g23849,g22771,g17868);
  and AND2_2550(g23851,g7329,g23048);
  and AND2_2551(g23852,g19179,g22696);
  and AND2_2552(g23854,g18265,g23049);
  and AND2_2553(g23855,g22954,g9767);
  and AND2_2554(g23857,g14263,g23056);
  and AND2_2555(g23859,g22958,g9787);
  and AND2_2556(g23860,g22962,g9790);
  and AND2_2557(g23864,g18297,g23057);
  and AND2_2558(g23865,g22966,g9816);
  and AND2_2559(g23866,g22971,g9819);
  and AND2_2560(g23877,g18314,g23060);
  and AND2_2561(g23878,g22975,g9880);
  and AND2_2562(g23886,g18341,g23064);
  and AND2_2563(g23888,g18358,g23069);
  and AND2_2564(g23889,g22962,g9913);
  and AND2_2565(g23891,g14385,g23074);
  and AND2_2566(g23893,g22966,g9933);
  and AND2_2567(g23894,g22971,g9936);
  and AND2_2568(g23898,g18390,g23075);
  and AND2_2569(g23899,g22975,g9962);
  and AND2_2570(g23900,g22980,g9965);
  and AND2_2571(g23904,g3010,g22750);
  and AND2_2572(g23907,g18436,g23079);
  and AND2_2573(g23909,g18453,g23082);
  and AND2_2574(g23910,g22971,g10067);
  and AND2_2575(g23912,g14497,g23087);
  and AND2_2576(g23914,g22975,g10087);
  and AND2_2577(g23915,g22980,g10090);
  and AND2_2578(g23917,g7545,g23088);
  and AND2_2579(g23939,g18509,g23095);
  and AND2_2580(g23941,g18526,g23098);
  and AND2_2581(g23942,g22980,g10176);
  and AND2_2582(g23944,g7570,g23103);
  and AND2_2583(g23971,g18573,g23112);
  and AND2_2584(g23972,g2903,g23115);
  and AND2_2585(g24029,g2900,g22903);
  and AND2_2586(g24211,g22014,g10969);
  and AND2_2587(g24217,g22825,g10999);
  and AND2_2588(g24221,g22979,g11042);
  and AND2_2589(g24224,g22219,g11045);
  and AND2_2590(g24229,g22232,g11105);
  and AND2_2591(g24236,g22243,g11157);
  and AND2_2592(g24241,g22259,g11228);
  and AND2_2593(g24246,g21982,g11291);
  and AND2_2594(g24247,g22551,g11297);
  and AND2_2595(g24253,g21995,g11370);
  and AND2_2596(g24256,g22003,g11438);
  and AND3_221(g24427,g17086,g24134,g13626);
  and AND2_2597(g24429,g24115,g13614);
  and AND3_222(g24431,g17124,g24153,g13637);
  and AND3_223(g24432,g14642,g15904,g24115);
  and AND2_2598(g24433,g24134,g13626);
  and AND3_224(g24435,g17151,g24168,g13649);
  and AND3_225(g24436,g14669,g15933,g24134);
  and AND2_2599(g24437,g24153,g13637);
  and AND3_226(g24439,g14703,g15962,g24153);
  and AND2_2600(g24440,g24168,g13649);
  and AND3_227(g24441,g14737,g15981,g24168);
  and AND3_228(g24478,g23545,g21119,g21227);
  and AND3_229(g24529,g19933,g17896,g23403);
  and AND3_230(g24540,g18548,g23089,g23403);
  and AND3_231(g24541,g23420,g17896,g23052);
  and AND3_232(g24542,g19950,g18007,g23410);
  and AND3_233(g24550,g18548,g23420,g19948);
  and AND3_234(g24552,g18598,g23107,g23410);
  and AND3_235(g24553,g23429,g18007,g23071);
  and AND3_236(g24554,g19977,g18124,g23415);
  and AND2_2601(g24559,g79,g23448);
  and AND3_237(g24561,g18598,g23429,g19975);
  and AND3_238(g24563,g18630,g23120,g23415);
  and AND3_239(g24564,g23435,g18124,g23084);
  and AND3_240(g24565,g20007,g18240,g23424);
  and AND2_2602(g24569,g767,g23455);
  and AND3_241(g24571,g18630,g23435,g20005);
  and AND3_242(g24573,g18639,g23129,g23424);
  and AND3_243(g24574,g23441,g18240,g23100);
  and AND2_2603(g24578,g1453,g23464);
  and AND3_244(g24580,g18639,g23441,g20043);
  and AND2_2604(g24585,g2147,g23473);
  and AND2_2605(g24590,g23486,g23478);
  and AND2_2606(g24591,g83,g23853);
  and AND2_2607(g24595,g23502,g23489);
  and AND2_2608(g24596,g771,g23887);
  and AND2_2609(g24603,g23518,g23505);
  and AND2_2610(g24604,g1457,g23908);
  and AND2_2611(g24610,g23533,g23521);
  and AND2_2612(g24611,g2151,g23940);
  and AND2_2613(g24644,g17203,g24115);
  and AND2_2614(g24664,g17208,g24134);
  and AND2_2615(g24676,g13568,g24115);
  and AND2_2616(g24683,g17214,g24153);
  and AND2_2617(g24695,g13576,g24134);
  and AND2_2618(g24700,g17217,g24168);
  and AND2_2619(g24712,g13585,g24153);
  and AND2_2620(g24723,g13605,g24168);
  and AND2_2621(g24745,g15454,g24096);
  and AND2_2622(g24746,g15454,g24098);
  and AND2_2623(g24747,g9427,g24099);
  and AND2_2624(g24748,g672,g24101);
  and AND2_2625(g24749,g15540,g24102);
  and AND2_2626(g24750,g15454,g24104);
  and AND2_2627(g24751,g9427,g24105);
  and AND2_2628(g24752,g9507,g24106);
  and AND2_2629(g24754,g15540,g24107);
  and AND2_2630(g24755,g9569,g24108);
  and AND2_2631(g24757,g1358,g24110);
  and AND2_2632(g24758,g15618,g24111);
  and AND2_2633(g24759,g21825,g23885);
  and AND2_2634(g24760,g9427,g24112);
  and AND2_2635(g24761,g9507,g24113);
  and AND2_2636(g24762,g12876,g24114);
  and AND2_2637(g24767,g15540,g24121);
  and AND2_2638(g24768,g9569,g24122);
  and AND2_2639(g24769,g9649,g24123);
  and AND2_2640(g24772,g15618,g24124);
  and AND2_2641(g24773,g9711,g24125);
  and AND2_2642(g24774,g2052,g24127);
  and AND2_2643(g24775,g15694,g24128);
  and AND2_2644(g24776,g9507,g24129);
  and AND2_2645(g24777,g12876,g24130);
  and AND2_2646(g24779,g9569,g24131);
  and AND2_2647(g24780,g9649,g24132);
  and AND2_2648(g24781,g12916,g24133);
  and AND2_2649(g24788,g15618,g24140);
  and AND2_2650(g24789,g9711,g24141);
  and AND2_2651(g24790,g9795,g24142);
  and AND2_2652(g24792,g15694,g24143);
  and AND2_2653(g24793,g9857,g24144);
  and AND2_2654(g24794,g2746,g24146);
  and AND2_2655(g24795,g12017,g24232);
  and AND2_2656(g24796,g12876,g24147);
  and AND2_2657(g24798,g9649,g24148);
  and AND2_2658(g24799,g12916,g24149);
  and AND2_2659(g24802,g9711,g24150);
  and AND2_2660(g24803,g9795,g24151);
  and AND2_2661(g24804,g12945,g24152);
  and AND2_2662(g24809,g15694,g24159);
  and AND2_2663(g24810,g9857,g24160);
  and AND2_2664(g24811,g9941,g24161);
  and AND2_2665(g24813,g21825,g23905);
  and AND2_2666(g24818,g12916,g24162);
  and AND2_2667(g24821,g9795,g24163);
  and AND2_2668(g24822,g12945,g24164);
  and AND2_2669(g24824,g9857,g24165);
  and AND2_2670(g24825,g9941,g24166);
  and AND2_2671(g24826,g12974,g24167);
  and AND2_2672(g24831,g24100,g20401);
  and AND2_2673(g24838,g12945,g24175);
  and AND2_2674(g24840,g9941,g24176);
  and AND2_2675(g24841,g12974,g24177);
  and AND2_2676(g24843,g21825,g23918);
  and AND2_2677(g24846,g24109,g20426);
  and AND2_2678(g24853,g12974,g24180);
  and AND2_2679(g24855,g18174,g23731);
  and AND2_2680(g24858,g24047,g18873);
  and AND2_2681(g24861,g24126,g20448);
  and AND2_2682(g24867,g666,g23779);
  and AND2_2683(g24869,g24047,g18894);
  and AND2_2684(g24870,g18281,g23786);
  and AND2_2685(g24874,g24060,g18899);
  and AND2_2686(g24876,g24145,g20467);
  and AND2_2687(g24878,g19830,g24210);
  and AND2_2688(g24881,g24047,g18912);
  and AND2_2689(g24882,g1352,g23832);
  and AND2_2690(g24884,g24060,g18917);
  and AND2_2691(g24885,g18374,g23839);
  and AND2_2692(g24888,g24073,g18922);
  and AND2_2693(g24898,g24060,g18931);
  and AND2_2694(g24899,g2046,g23867);
  and AND2_2695(g24901,g24073,g18936);
  and AND2_2696(g24902,g18469,g23874);
  and AND2_2697(g24905,g24084,g18941);
  and AND2_2698(g24906,g18886,g23879);
  and AND2_2699(g24907,g7466,g24220);
  and AND2_2700(g24908,g7342,g23882);
  and AND2_2701(g24921,g24073,g18951);
  and AND2_2702(g24922,g2740,g23901);
  and AND2_2703(g24924,g24084,g18956);
  and AND2_2704(g24938,g24084,g18967);
  and AND2_2705(g24964,g7595,g24251);
  and AND2_2706(g24974,g7600,g24030);
  and AND2_2707(g25086,g23444,g10880);
  and AND2_2708(g25102,g23444,g10915);
  and AND2_2709(g25117,g23444,g10974);
  and AND3_245(g25128,g17051,g24115,g13614);
  and AND2_2710(g25178,g24623,g20634);
  and AND2_2711(g25181,g24636,g20673);
  and AND2_2712(g25182,g24681,g20676);
  and AND2_2713(g25184,g24694,g20735);
  and AND2_2714(g25187,g24633,g16608);
  and AND2_2715(g25188,g24652,g20763);
  and AND2_2716(g25192,g24711,g20790);
  and AND2_2717(g25193,g24653,g16626);
  and AND2_2718(g25196,g24672,g16640);
  and AND2_2719(g25198,g24691,g16651);
  and AND2_2720(g25269,g24648,g8700);
  and AND2_2721(g25277,g24648,g8714);
  and AND2_2722(g25278,g24668,g8719);
  and AND2_2723(g25281,g5606,g24815);
  and AND2_2724(g25282,g24648,g8748);
  and AND2_2725(g25286,g24668,g8752);
  and AND2_2726(g25287,g24687,g8757);
  and AND2_2727(g25289,g5631,g24834);
  and AND2_2728(g25290,g24668,g8771);
  and AND2_2729(g25294,g24687,g8775);
  and AND2_2730(g25295,g24704,g8780);
  and AND2_2731(g25299,g5659,g24850);
  and AND2_2732(g25300,g24687,g8794);
  and AND2_2733(g25304,g24704,g8798);
  and AND2_2734(g25309,g5697,g24864);
  and AND2_2735(g25310,g24704,g8813);
  and AND3_246(g25318,g24682,g19358,g19335);
  and AND2_2736(g25321,g25075,g9669);
  and AND2_2737(g25328,g24644,g17892);
  and AND2_2738(g25334,g24644,g17984);
  and AND2_2739(g25337,g24664,g18003);
  and AND2_2740(g25342,g5851,g24600);
  and AND2_2741(g25346,g24644,g18084);
  and AND2_2742(g25348,g24664,g18101);
  and AND2_2743(g25351,g24683,g18120);
  and AND2_2744(g25356,g5898,g24607);
  and AND2_2745(g25360,g24664,g18200);
  and AND2_2746(g25362,g24683,g18217);
  and AND2_2747(g25365,g24700,g18236);
  and AND2_2748(g25371,g5937,g24619);
  and AND2_2749(g25375,g24683,g18307);
  and AND2_2750(g25377,g24700,g18324);
  and AND2_2751(g25388,g5971,g24630);
  and AND2_2752(g25392,g24700,g18400);
  and AND2_2753(g25453,g6142,g24763);
  and AND2_2754(g25457,g6163,g24784);
  and AND2_2755(g25461,g6190,g24805);
  and AND2_2756(g25466,g6222,g24827);
  and AND2_2757(g25470,g24479,g20400);
  and AND2_2758(g25475,g14148,g25087);
  and AND2_2759(g25482,g24480,g17567);
  and AND2_2760(g25483,g24481,g20421);
  and AND2_2761(g25487,g24485,g20425);
  and AND2_2762(g25505,g6707,g25094);
  and AND2_2763(g25506,g14263,g25095);
  and AND2_2764(g25513,g24487,g17664);
  and AND2_2765(g25514,g24488,g20443);
  and AND2_2766(g25518,g24489,g20447);
  and AND2_2767(g25552,g7009,g25104);
  and AND2_2768(g25553,g14385,g25105);
  and AND2_2769(g25560,g24494,g17764);
  and AND2_2770(g25561,g24495,g20462);
  and AND2_2771(g25565,g24496,g20466);
  and AND2_2772(g25618,g7259,g25110);
  and AND2_2773(g25619,g14497,g25111);
  and AND2_2774(g25626,g24504,g17865);
  and AND2_2775(g25627,g24505,g20477);
  and AND2_2776(g25628,g21008,g25115);
  and AND2_2777(g25629,g3024,g25116);
  and AND2_2778(g25697,g7455,g25120);
  and AND2_2779(g25881,g2908,g25126);
  and AND2_2780(g25951,g24800,g13670);
  and AND2_2781(g25953,g24783,g13699);
  and AND2_2782(g25957,g24782,g11869);
  and AND2_2783(g25961,g24770,g11901);
  and AND2_2784(g25963,g24756,g11944);
  and AND2_2785(g25968,g24871,g11986);
  and AND2_2786(g25972,g24859,g12042);
  and AND2_2787(g25973,g24847,g13838);
  and AND2_2788(g25975,g24606,g21917);
  and AND2_2789(g25977,g24845,g12089);
  and AND2_2790(g25978,g24836,g13850);
  and AND2_2791(g25980,g24663,g21928);
  and AND2_2792(g25981,g24819,g13858);
  and AND2_2793(g26023,g25422,g24912);
  and AND2_2794(g26024,g25301,g21102);
  and AND2_2795(g26026,g25431,g24929);
  and AND2_2796(g26027,g25418,g22271);
  and AND2_2797(g26028,g25438,g24941);
  and AND2_2798(g26029,g25445,g24952);
  and AND2_2799(g26030,g25429,g22304);
  and AND2_2800(g26032,g25379,g19415);
  and AND2_2801(g26033,g25395,g19452);
  and AND2_2802(g26034,g25405,g19479);
  and AND2_2803(g26035,g25523,g19483);
  and AND2_2804(g26036,g25413,g19502);
  and AND2_2805(g26038,g25589,g19504);
  and AND2_2806(g26039,g25668,g19523);
  and AND2_2807(g26040,g25745,g19533);
  and AND2_2808(g26051,g70,g25296);
  and AND2_2809(g26052,g25941,g21087);
  and AND2_2810(g26053,g758,g25306);
  and AND2_2811(g26054,g25944,g21099);
  and AND2_2812(g26060,g25943,g21108);
  and AND2_2813(g26061,g1444,g25315);
  and AND2_2814(g26062,g25947,g21113);
  and AND2_2815(g26067,g25946,g21125);
  and AND2_2816(g26068,g2138,g25324);
  and AND2_2817(g26069,g25949,g21130);
  and AND2_2818(g26074,g25948,g21144);
  and AND2_2819(g26075,g74,g25698);
  and AND2_2820(g26080,g25950,g21164);
  and AND2_2821(g26082,g762,g25771);
  and AND2_2822(g26085,g1448,g25825);
  and AND2_2823(g26091,g2142,g25860);
  and AND2_2824(g26157,g21825,g25630);
  and AND2_2825(g26158,g679,g25937);
  and AND2_2826(g26163,g1365,g25939);
  and AND2_2827(g26166,g686,g25454);
  and AND2_2828(g26171,g2059,g25942);
  and AND2_2829(g26186,g1372,g25458);
  and AND2_2830(g26188,g2753,g25945);
  and AND2_2831(g26207,g2066,g25463);
  and AND2_2832(g26212,g4217,g25467);
  and AND2_2833(g26213,g25895,g9306);
  and AND2_2834(g26231,g2760,g25472);
  and AND2_2835(g26233,g4340,g25476);
  and AND2_2836(g26234,g4343,g25479);
  and AND2_2837(g26235,g25895,g9368);
  and AND2_2838(g26236,g25899,g9371);
  and AND2_2839(g26243,g4372,g25484);
  and AND2_2840(g26244,g25903,g9387);
  and AND2_2841(g26257,g4465,g25493);
  and AND2_2842(g26258,g4468,g25496);
  and AND2_2843(g26259,g4471,g25499);
  and AND2_2844(g26260,g25254,g17649);
  and AND2_2845(g26261,g25895,g9443);
  and AND2_2846(g26262,g25899,g9446);
  and AND2_2847(g26263,g4476,g25502);
  and AND2_2848(g26268,g4509,g25507);
  and AND2_2849(g26269,g4512,g25510);
  and AND2_2850(g26270,g25903,g9465);
  and AND2_2851(g26271,g25907,g9468);
  and AND2_2852(g26278,g4541,g25515);
  and AND2_2853(g26279,g25911,g9484);
  and AND2_2854(g26288,g4592,g25524);
  and AND2_2855(g26289,g4595,g25527);
  and AND2_2856(g26290,g4598,g25530);
  and AND2_2857(g26291,g25899,g9524);
  and AND2_2858(g26292,g4603,g25533);
  and AND2_2859(g26293,g4606,g25536);
  and AND2_2860(g26298,g4641,g25540);
  and AND2_2861(g26299,g4644,g25543);
  and AND2_2862(g26300,g4647,g25546);
  and AND2_2863(g26301,g25258,g17749);
  and AND2_2864(g26302,g25903,g9585);
  and AND2_2865(g26303,g25907,g9588);
  and AND2_2866(g26307,g4652,g25549);
  and AND2_2867(g26309,g4685,g25554);
  and AND2_2868(g26310,g4688,g25557);
  and AND2_2869(g26311,g25911,g9607);
  and AND2_2870(g26312,g25915,g9610);
  and AND2_2871(g26316,g4717,g25562);
  and AND2_2872(g26317,g25919,g9626);
  and AND2_2873(g26318,g4737,g25573);
  and AND2_2874(g26319,g4740,g25576);
  and AND2_2875(g26324,g4743,g25579);
  and AND2_2876(g26325,g4746,g25582);
  and AND2_2877(g26326,g4749,g25585);
  and AND2_2878(g26332,g4769,g25590);
  and AND2_2879(g26333,g4772,g25593);
  and AND2_2880(g26334,g4775,g25596);
  and AND2_2881(g26335,g25907,g9666);
  and AND2_2882(g26339,g4780,g25599);
  and AND2_2883(g26340,g4783,g25602);
  and AND2_2884(g26342,g4818,g25606);
  and AND2_2885(g26343,g4821,g25609);
  and AND2_2886(g26344,g4824,g25612);
  and AND2_2887(g26345,g25261,g17850);
  and AND2_2888(g26346,g25911,g9727);
  and AND2_2889(g26347,g25915,g9730);
  and AND2_2890(g26348,g4829,g25615);
  and AND2_2891(g26350,g4862,g25620);
  and AND2_2892(g26351,g4865,g25623);
  and AND2_2893(g26352,g25919,g9749);
  and AND2_2894(g26353,g25923,g9752);
  and AND2_2895(g26357,g4882,g25634);
  and AND2_2896(g26361,g4888,g25637);
  and AND2_2897(g26362,g4891,g25640);
  and AND2_2898(g26363,g4894,g25643);
  and AND2_2899(g26365,g4913,g25652);
  and AND2_2900(g26366,g4916,g25655);
  and AND2_2901(g26371,g4919,g25658);
  and AND2_2902(g26372,g4922,g25661);
  and AND2_2903(g26373,g4925,g25664);
  and AND2_2904(g26379,g4945,g25669);
  and AND2_2905(g26380,g4948,g25672);
  and AND2_2906(g26381,g4951,g25675);
  and AND2_2907(g26382,g25915,g9812);
  and AND2_2908(g26383,g4956,g25678);
  and AND2_2909(g26384,g4959,g25681);
  and AND2_2910(g26386,g4994,g25685);
  and AND2_2911(g26387,g4997,g25688);
  and AND2_2912(g26388,g5000,g25691);
  and AND2_2913(g26389,g25264,g17962);
  and AND2_2914(g26390,g25919,g9873);
  and AND2_2915(g26391,g25923,g9876);
  and AND2_2916(g26392,g5005,g25694);
  and AND2_2917(g26396,g5027,g25700);
  and AND2_2918(g26397,g5030,g25703);
  and AND2_2919(g26400,g5041,g25711);
  and AND2_2920(g26404,g5047,g25714);
  and AND2_2921(g26405,g5050,g25717);
  and AND2_2922(g26406,g5053,g25720);
  and AND2_2923(g26408,g5072,g25729);
  and AND2_2924(g26409,g5075,g25732);
  and AND2_2925(g26414,g5078,g25735);
  and AND2_2926(g26415,g5081,g25738);
  and AND2_2927(g26416,g5084,g25741);
  and AND2_2928(g26422,g5104,g25746);
  and AND2_2929(g26423,g5107,g25749);
  and AND2_2930(g26424,g5110,g25752);
  and AND2_2931(g26425,g25923,g9958);
  and AND2_2932(g26426,g5115,g25755);
  and AND2_2933(g26427,g5118,g25758);
  and AND2_2934(g26432,g5145,g25767);
  and AND2_2935(g26437,g5156,g25773);
  and AND2_2936(g26438,g5159,g25776);
  and AND2_2937(g26441,g5170,g25784);
  and AND2_2938(g26445,g5176,g25787);
  and AND2_2939(g26446,g5179,g25790);
  and AND2_2940(g26447,g5182,g25793);
  and AND2_2941(g26449,g5201,g25802);
  and AND2_2942(g26450,g5204,g25805);
  and AND2_2943(g26455,g5207,g25808);
  and AND2_2944(g26456,g5210,g25811);
  and AND2_2945(g26457,g5213,g25814);
  and AND2_2946(g26464,g5238,g25821);
  and AND2_2947(g26469,g5249,g25827);
  and AND2_2948(g26470,g5252,g25830);
  and AND2_2949(g26473,g5263,g25838);
  and AND2_2950(g26477,g5269,g25841);
  and AND2_2951(g26478,g5272,g25844);
  and AND2_2952(g26479,g5275,g25847);
  and AND2_2953(g26488,g5301,g25856);
  and AND2_2954(g26493,g5312,g25862);
  and AND2_2955(g26494,g5315,g25865);
  and AND2_2956(g26504,g5338,g25877);
  and AND2_2957(g26663,g25274,g21066);
  and AND2_2958(g26668,g25283,g21076);
  and AND2_2959(g26673,g12431,g25318);
  and AND2_2960(g26674,g25291,g21090);
  and AND2_2961(g26754,g14657,g26508);
  and AND2_2962(g26755,g26083,g22239);
  and AND2_2963(g26756,g26113,g22240);
  and AND3_247(g26758,g16614,g26521,g13637);
  and AND2_2964(g26759,g26356,g19251);
  and AND2_2965(g26760,g26137,g22256);
  and AND2_2966(g26761,g26154,g22257);
  and AND2_2967(g26763,g14691,g26516);
  and AND3_248(g26764,g16632,g26525,g13649);
  and AND2_2968(g26765,g26399,g19265);
  and AND2_2969(g26766,g14725,g26521);
  and AND2_2970(g26767,g26087,g22287);
  and AND2_2971(g26768,g26440,g19280);
  and AND2_2972(g26769,g14753,g26525);
  and AND2_2973(g26770,g26059,g19287);
  and AND3_249(g26771,g24912,g26508,g13614);
  and AND2_2974(g26773,g26145,g22303);
  and AND2_2975(g26774,g26472,g19299);
  and AND2_2976(g26775,g26099,g22318);
  and AND2_2977(g26777,g26066,g19305);
  and AND3_250(g26778,g24929,g26516,g13626);
  and AND2_2978(g26780,g26119,g16622);
  and AND2_2979(g26783,g26073,g19326);
  and AND3_251(g26784,g24941,g26521,g13637);
  and AND2_2980(g26787,g26129,g16636);
  and AND2_2981(g26790,g26079,g19353);
  and AND3_252(g26791,g24952,g26525,g13649);
  and AND2_2982(g26794,g26143,g16647);
  and AND2_2983(g26797,g26148,g16659);
  and AND2_2984(g26829,g5623,g26209);
  and AND2_2985(g26833,g5651,g26237);
  and AND2_2986(g26842,g5689,g26275);
  and AND2_2987(g26845,g5664,g26056);
  and AND2_2988(g26851,g5741,g26313);
  and AND2_2989(g26853,g5716,g26063);
  and AND2_2990(g26860,g5774,g26070);
  and AND2_2991(g26866,g5833,g26076);
  and AND2_2992(g26955,g6157,g26533);
  and AND2_2993(g26958,g6184,g26538);
  and AND2_2994(g26961,g13907,g26175);
  and AND2_2995(g26962,g6180,g26178);
  and AND2_2996(g26963,g6216,g26539);
  and AND2_2997(g26965,g23320,g26540);
  and AND2_2998(g26966,g13963,g26196);
  and AND2_2999(g26967,g6212,g26202);
  and AND2_3000(g26968,g6305,g26542);
  and AND2_3001(g26969,g23320,g26543);
  and AND2_3002(g26970,g21976,g26544);
  and AND2_3003(g26971,g23325,g26546);
  and AND2_3004(g26972,g14033,g26223);
  and AND2_3005(g26973,g6301,g26226);
  and AND2_3006(g26977,g23320,g26550);
  and AND2_3007(g26978,g21976,g26551);
  and AND2_3008(g26979,g23331,g26552);
  and AND2_3009(g26980,g23360,g26554);
  and AND2_3010(g26981,g23325,g26555);
  and AND2_3011(g26982,g21983,g26556);
  and AND2_3012(g26984,g23335,g26558);
  and AND2_3013(g26985,g14124,g26251);
  and AND2_3014(g26986,g6438,g26254);
  and AND2_3015(g26993,g21976,g26561);
  and AND2_3016(g26994,g23331,g26562);
  and AND2_3017(g26995,g21991,g26563);
  and AND2_3018(g26996,g23360,g26564);
  and AND2_3019(g26997,g22050,g26565);
  and AND2_3020(g26998,g23325,g26566);
  and AND2_3021(g26999,g21983,g26567);
  and AND2_3022(g27000,g23340,g26568);
  and AND2_3023(g27001,g23364,g26570);
  and AND2_3024(g27002,g23335,g26571);
  and AND2_3025(g27003,g21996,g26572);
  and AND2_3026(g27004,g23344,g26574);
  and AND2_3027(g27005,g23331,g26578);
  and AND2_3028(g27006,g21991,g26579);
  and AND2_3029(g27007,g23360,g26580);
  and AND2_3030(g27008,g22050,g26581);
  and AND2_3031(g27009,g23368,g26582);
  and AND2_3032(g27016,g21983,g26584);
  and AND2_3033(g27017,g23340,g26585);
  and AND2_3034(g27018,g22005,g26586);
  and AND2_3035(g27019,g23364,g26587);
  and AND2_3036(g27020,g22069,g26588);
  and AND2_3037(g27021,g23335,g26589);
  and AND2_3038(g27022,g21996,g26590);
  and AND2_3039(g27023,g23349,g26591);
  and AND2_3040(g27024,g23372,g26593);
  and AND2_3041(g27025,g23344,g26594);
  and AND2_3042(g27026,g22009,g26595);
  and AND2_3043(g27027,g21991,g26598);
  and AND2_3044(g27028,g22050,g26599);
  and AND2_3045(g27029,g23368,g26600);
  and AND2_3046(g27030,g22083,g26601);
  and AND2_3047(g27031,g23340,g26602);
  and AND2_3048(g27032,g22005,g26603);
  and AND2_3049(g27033,g23364,g26604);
  and AND2_3050(g27034,g22069,g26605);
  and AND2_3051(g27035,g23377,g26606);
  and AND2_3052(g27042,g21996,g26608);
  and AND2_3053(g27043,g23349,g26609);
  and AND2_3054(g27044,g22016,g26610);
  and AND2_3055(g27045,g23372,g26611);
  and AND2_3056(g27046,g22093,g26612);
  and AND2_3057(g27047,g23344,g26613);
  and AND2_3058(g27048,g22009,g26614);
  and AND2_3059(g27049,g23353,g26615);
  and AND2_3060(g27050,g23381,g26617);
  and AND2_3061(g27052,g4885,g26358);
  and AND2_3062(g27053,g23368,g26619);
  and AND2_3063(g27054,g22083,g26620);
  and AND2_3064(g27055,g22005,g26621);
  and AND2_3065(g27056,g22069,g26622);
  and AND2_3066(g27057,g23377,g26623);
  and AND2_3067(g27058,g22108,g26624);
  and AND2_3068(g27059,g23349,g26625);
  and AND2_3069(g27060,g22016,g26626);
  and AND2_3070(g27061,g23372,g26627);
  and AND2_3071(g27062,g22093,g26628);
  and AND2_3072(g27063,g23388,g26629);
  and AND2_3073(g27070,g22009,g26631);
  and AND2_3074(g27071,g23353,g26632);
  and AND2_3075(g27072,g22021,g26633);
  and AND2_3076(g27073,g23381,g26634);
  and AND2_3077(g27074,g22118,g26635);
  and AND2_3078(g27076,g5024,g26393);
  and AND2_3079(g27077,g22083,g26636);
  and AND2_3080(g27079,g5044,g26401);
  and AND2_3081(g27080,g23377,g26637);
  and AND2_3082(g27081,g22108,g26638);
  and AND2_3083(g27082,g22016,g26639);
  and AND2_3084(g27083,g22093,g26640);
  and AND2_3085(g27084,g23388,g26641);
  and AND2_3086(g27085,g22134,g26642);
  and AND2_3087(g27086,g23353,g26643);
  and AND2_3088(g27087,g22021,g26644);
  and AND2_3089(g27088,g23381,g26645);
  and AND2_3090(g27089,g22118,g26646);
  and AND2_3091(g27090,g23395,g26647);
  and AND2_3092(g27091,g5142,g26429);
  and AND2_3093(g27092,g5153,g26434);
  and AND2_3094(g27093,g22108,g26648);
  and AND2_3095(g27095,g5173,g26442);
  and AND2_3096(g27096,g23388,g26649);
  and AND2_3097(g27097,g22134,g26650);
  and AND2_3098(g27098,g22021,g26651);
  and AND2_3099(g27099,g22118,g26652);
  and AND2_3100(g27100,g23395,g26653);
  and AND2_3101(g27101,g22157,g26654);
  and AND2_3102(g27103,g5235,g26461);
  and AND2_3103(g27104,g5246,g26466);
  and AND2_3104(g27105,g22134,g26656);
  and AND2_3105(g27107,g5266,g26474);
  and AND2_3106(g27108,g23395,g26657);
  and AND2_3107(g27109,g22157,g26658);
  and AND2_3108(g27110,g5298,g26485);
  and AND2_3109(g27111,g5309,g26490);
  and AND2_3110(g27112,g22157,g26662);
  and AND2_3111(g27115,g5335,g26501);
  and AND2_3112(g27178,g26110,g22213);
  and AND3_253(g27181,g16570,g26508,g13614);
  and AND2_3113(g27182,g26151,g22217);
  and AND2_3114(g27185,g26126,g22230);
  and AND3_254(g27187,g16594,g26516,g13626);
  and AND2_3115(g27240,g26905,g22241);
  and AND2_3116(g27241,g10730,g26934);
  and AND2_3117(g27242,g26793,g8357);
  and AND2_3118(g27244,g26914,g22258);
  and AND2_3119(g27245,g26877,g22286);
  and AND2_3120(g27246,g26988,g16676);
  and AND2_3121(g27247,g27011,g16702);
  and AND2_3122(g27248,g27037,g16733);
  and AND2_3123(g27249,g27065,g16775);
  and AND2_3124(g27355,g61,g26837);
  and AND2_3125(g27356,g65,g26987);
  and AND2_3126(g27358,g749,g26846);
  and AND2_3127(g27359,g753,g27010);
  and AND2_3128(g27364,g1435,g26855);
  and AND2_3129(g27365,g1439,g27036);
  and AND2_3130(g27370,g27126,g8874);
  and AND2_3131(g27371,g2129,g26861);
  and AND2_3132(g27372,g2133,g27064);
  and AND2_3133(g27394,g17802,g27134);
  and AND2_3134(g27396,g692,g27135);
  and AND2_3135(g27407,g17914,g27136);
  and AND2_3136(g27409,g1378,g27137);
  and AND2_3137(g27425,g18025,g27138);
  and AND2_3138(g27427,g2072,g27139);
  and AND2_3139(g27446,g18142,g27141);
  and AND2_3140(g27448,g2766,g27142);
  and AND2_3141(g27495,g23945,g27146);
  and AND2_3142(g27509,g23945,g27148);
  and AND2_3143(g27516,g23974,g27151);
  and AND2_3144(g27530,g23945,g27153);
  and AND2_3145(g27534,g23974,g27155);
  and AND2_3146(g27541,g24004,g27159);
  and AND2_3147(g27552,g23974,g27162);
  and AND2_3148(g27554,g24004,g27164);
  and AND2_3149(g27561,g24038,g27167);
  and AND2_3150(g27568,g24004,g27172);
  and AND2_3151(g27570,g24038,g27173);
  and AND2_3152(g27578,g24038,g27177);
  and AND2_3153(g27656,g26796,g11004);
  and AND2_3154(g27657,g27114,g11051);
  and AND2_3155(g27659,g27132,g11114);
  and AND2_3156(g27660,g26835,g11117);
  and AND2_3157(g27661,g26841,g11173);
  and AND2_3158(g27666,g26849,g11243);
  and AND2_3159(g27671,g26885,g22212);
  and AND2_3160(g27673,g26854,g11312);
  and AND2_3161(g27679,g26782,g11386);
  and AND2_3162(g27680,g26983,g11392);
  and AND2_3163(g27681,g26788,g11456);
  and AND2_3164(g27719,g27496,g20649);
  and AND2_3165(g27720,g27481,g20652);
  and AND2_3166(g27721,g27579,g20655);
  and AND2_3167(g27723,g27464,g20679);
  and AND2_3168(g27725,g27532,g20704);
  and AND2_3169(g27726,g27531,g20732);
  and AND2_3170(g27727,g27414,g19301);
  and AND2_3171(g27728,g27564,g20766);
  and AND2_3172(g27729,g27435,g19322);
  and AND2_3173(g27730,g27454,g19349);
  and AND2_3174(g27731,g27470,g19383);
  and AND2_3175(g27732,g27492,g16758);
  and AND2_3176(g27733,g27513,g16785);
  and AND2_3177(g27734,g27538,g16814);
  and AND2_3178(g27737,g27558,g16832);
  and AND2_3179(g27770,g5642,g27449);
  and AND2_3180(g27772,g5680,g27465);
  and AND2_3181(g27773,g5732,g27484);
  and AND2_3182(g27774,g5702,g27361);
  and AND2_3183(g27775,g5790,g27506);
  and AND2_3184(g27779,g5760,g27367);
  and AND2_3185(g27783,g5819,g27373);
  and AND2_3186(g27790,g5875,g27376);
  and AND2_3187(g27904,g13873,g27387);
  and AND2_3188(g27908,g13886,g27391);
  and AND2_3189(g27909,g13895,g27397);
  and AND2_3190(g27913,g4017,g27401);
  and AND2_3191(g27914,g13927,g27404);
  and AND2_3192(g27915,g13936,g27410);
  and AND2_3193(g27922,g4112,g27416);
  and AND2_3194(g27923,g4144,g27419);
  and AND2_3195(g27924,g13983,g27422);
  and AND2_3196(g27926,g13992,g27428);
  and AND2_3197(g27931,g4221,g27432);
  and AND2_3198(g27935,g4251,g27437);
  and AND2_3199(g27936,g4283,g27440);
  and AND2_3200(g27938,g14053,g27443);
  and AND2_3201(g27945,g4376,g27451);
  and AND2_3202(g27949,g4406,g27456);
  and AND2_3203(g27951,g4438,g27459);
  and AND2_3204(g27963,g4545,g27467);
  and AND2_3205(g27968,g4575,g27472);
  and AND2_3206(g27970,g14238,g27475);
  and AND2_3207(g27984,g4721,g27486);
  and AND2_3208(g27985,g14342,g27489);
  and AND2_3209(g27991,g14360,g27498);
  and AND2_3210(g28008,g27590,g9770);
  and AND2_3211(g28009,g14454,g27510);
  and AND2_3212(g28015,g14472,g27518);
  and AND2_3213(g28027,g27590,g9895);
  and AND2_3214(g28028,g27595,g9898);
  and AND2_3215(g28035,g27599,g9916);
  and AND2_3216(g28036,g14541,g27535);
  and AND2_3217(g28042,g14559,g27543);
  and AND2_3218(g28050,g27590,g10018);
  and AND2_3219(g28051,g27595,g10021);
  and AND2_3220(g28057,g27599,g10049);
  and AND2_3221(g28058,g27604,g10052);
  and AND2_3222(g28065,g27608,g10070);
  and AND2_3223(g28066,g14596,g27555);
  and AND2_3224(g28073,g27595,g10109);
  and AND2_3225(g28079,g27599,g10127);
  and AND2_3226(g28080,g27604,g10130);
  and AND2_3227(g28086,g27608,g10158);
  and AND2_3228(g28087,g27613,g10161);
  and AND2_3229(g28094,g27617,g10179);
  and AND2_3230(g28098,g27604,g10214);
  and AND2_3231(g28104,g27608,g10232);
  and AND2_3232(g28105,g27613,g10235);
  and AND2_3233(g28111,g27617,g10263);
  and AND2_3234(g28112,g27622,g10266);
  and AND2_3235(g28116,g27613,g10316);
  and AND2_3236(g28122,g27617,g10334);
  and AND2_3237(g28123,g27622,g10337);
  and AND2_3238(g28127,g27622,g10409);
  and AND2_3239(g28171,g27349,g10898);
  and AND2_3240(g28176,g27349,g10940);
  and AND2_3241(g28188,g27349,g11008);
  and AND2_3242(g28193,g27573,g21914);
  and AND2_3243(g28319,g27855,g22246);
  and AND2_3244(g28320,g27854,g20637);
  and AND2_3245(g28322,g27937,g13868);
  and AND2_3246(g28323,g8580,g27838);
  and AND2_3247(g28324,g27810,g20659);
  and AND2_3248(g28326,g27865,g22274);
  and AND2_3249(g28327,g27900,g22275);
  and AND2_3250(g28329,g27823,g20708);
  and AND2_3251(g28330,g27864,g20711);
  and AND2_3252(g28331,g27802,g22307);
  and AND2_3253(g28332,g27883,g22331);
  and AND2_3254(g28333,g27882,g20772);
  and AND2_3255(g28334,g27842,g20793);
  and AND2_3256(g28335,g27814,g22343);
  and AND2_3257(g28336,g27896,g20810);
  and AND2_3258(g28337,g28002,g19448);
  and AND2_3259(g28338,g28029,g19475);
  and AND2_3260(g28339,g28059,g19498);
  and AND2_3261(g28340,g28088,g19519);
  and AND2_3262(g28373,g56,g27969);
  and AND2_3263(g28376,g744,g27990);
  and AND2_3264(g28378,g52,g27776);
  and AND3_255(g28379,g27868,g19390,g19369);
  and AND2_3265(g28380,g1430,g28014);
  and AND2_3266(g28381,g28157,g9815);
  and AND2_3267(g28383,g740,g27780);
  and AND2_3268(g28385,g2124,g28041);
  and AND2_3269(g28387,g1426,g27787);
  and AND2_3270(g28389,g2120,g27794);
  and AND2_3271(g28396,g7754,g27806);
  and AND2_3272(g28398,g7769,g27817);
  and AND2_3273(g28399,g7776,g27820);
  and AND2_3274(g28401,g7782,g27831);
  and AND2_3275(g28402,g7785,g27839);
  and AND2_3276(g28404,g7792,g27843);
  and AND2_3277(g28405,g7796,g27847);
  and AND2_3278(g28407,g7799,g27858);
  and AND2_3279(g28408,g7806,g27861);
  and AND2_3280(g28411,g7809,g27872);
  and AND2_3281(g28412,g7812,g27879);
  and AND2_3282(g28416,g7823,g27889);
  and AND2_3283(g28422,g17640,g28150);
  and AND2_3284(g28423,g17724,g28152);
  and AND2_3285(g28424,g17741,g28153);
  and AND2_3286(g28426,g28128,g9170);
  and AND2_3287(g28427,g26092,g28154);
  and AND2_3288(g28428,g17825,g28155);
  and AND2_3289(g28429,g17842,g28156);
  and AND2_3290(g28430,g28128,g9196);
  and AND2_3291(g28431,g26092,g28158);
  and AND2_3292(g28433,g28133,g9212);
  and AND2_3293(g28434,g26114,g28159);
  and AND2_3294(g28435,g17937,g28160);
  and AND2_3295(g28436,g17954,g28161);
  and AND2_3296(g28438,g17882,g27919);
  and AND2_3297(g28439,g28128,g9242);
  and AND2_3298(g28440,g26092,g28162);
  and AND2_3299(g28441,g28133,g9257);
  and AND2_3300(g28442,g26114,g28163);
  and AND2_3301(g28444,g28137,g9273);
  and AND2_3302(g28445,g26121,g28164);
  and AND2_3303(g28446,g18048,g28165);
  and AND2_3304(g28448,g17974,g27928);
  and AND2_3305(g28450,g17993,g27932);
  and AND2_3306(g28451,g28133,g9320);
  and AND2_3307(g28452,g26114,g28166);
  and AND2_3308(g28453,g28137,g9335);
  and AND2_3309(g28454,g26121,g28167);
  and AND2_3310(g28456,g28141,g9351);
  and AND2_3311(g28457,g26131,g28168);
  and AND2_3312(g28459,g18074,g27939);
  and AND2_3313(g28460,g18091,g27942);
  and AND2_3314(g28462,g18110,g27946);
  and AND2_3315(g28463,g28137,g9401);
  and AND2_3316(g28464,g26121,g28169);
  and AND2_3317(g28465,g28141,g9416);
  and AND2_3318(g28466,g26131,g28170);
  and AND2_3319(g28468,g18265,g28172);
  and AND2_3320(g28469,g18179,g27952);
  and AND2_3321(g28471,g18190,g27956);
  and AND2_3322(g28472,g18207,g27959);
  and AND2_3323(g28474,g18226,g27965);
  and AND2_3324(g28475,g28141,g9498);
  and AND2_3325(g28476,g26131,g28173);
  and AND2_3326(g28477,g18341,g28174);
  and AND2_3327(g28478,g18358,g28175);
  and AND2_3328(g28479,g18286,g27973);
  and AND2_3329(g28480,g18297,g27977);
  and AND2_3330(g28481,g18314,g27981);
  and AND2_3331(g28484,g18436,g28177);
  and AND2_3332(g28485,g18453,g28178);
  and AND2_3333(g28486,g18379,g27994);
  and AND2_3334(g28487,g18390,g27999);
  and AND2_3335(g28492,g18509,g28186);
  and AND2_3336(g28493,g18526,g28187);
  and AND2_3337(g28494,g18474,g28018);
  and AND2_3338(g28497,g18573,g28190);
  and AND2_3339(g28657,g27925,g13700);
  and AND2_3340(g28659,g27917,g13736);
  and AND2_3341(g28660,g27916,g11911);
  and AND2_3342(g28662,g27911,g11951);
  and AND2_3343(g28663,g27906,g11997);
  and AND2_3344(g28664,g27997,g12055);
  and AND2_3345(g28665,g27827,g22222);
  and AND2_3346(g28666,g27980,g12106);
  and AND2_3347(g28667,g27964,g13852);
  and AND2_3348(g28669,g27897,g22233);
  and AND2_3349(g28670,g27798,g21935);
  and AND2_3350(g28671,g27962,g12161);
  and AND2_3351(g28672,g27950,g13859);
  and AND2_3352(g28707,g12436,g28379);
  and AND2_3353(g28708,g28392,g22260);
  and AND2_3354(g28709,g28400,g22261);
  and AND2_3355(g28710,g28403,g22262);
  and AND2_3356(g28711,g10749,g28415);
  and AND2_3357(g28712,g28406,g22276);
  and AND2_3358(g28713,g28410,g22290);
  and AND2_3359(g28714,g28394,g22306);
  and AND2_3360(g28715,g28414,g22332);
  and AND2_3361(g28716,g28449,g19319);
  and AND2_3362(g28717,g28461,g19346);
  and AND2_3363(g28718,g28473,g19380);
  and AND2_3364(g28719,g28482,g19412);
  and AND2_3365(g28722,g28523,g16694);
  and AND2_3366(g28724,g28551,g16725);
  and AND2_3367(g28726,g28578,g16767);
  and AND2_3368(g28729,g28606,g16794);
  and AND2_3369(g28834,g5751,g28483);
  and AND2_3370(g28836,g5810,g28491);
  and AND2_3371(g28838,g5866,g28496);
  and AND2_3372(g28840,g5913,g28500);
  and AND2_3373(g28841,g27834,g28554);
  and AND2_3374(g28843,g27834,g28581);
  and AND2_3375(g28844,g27850,g28582);
  and AND2_3376(g28846,g27834,g28608);
  and AND2_3377(g28847,g27850,g28609);
  and AND2_3378(g28848,g27875,g28610);
  and AND2_3379(g28849,g27850,g28616);
  and AND2_3380(g28850,g27875,g28617);
  and AND2_3381(g28851,g27892,g28618);
  and AND2_3382(g28852,g27875,g28623);
  and AND2_3383(g28853,g27892,g28624);
  and AND2_3384(g28854,g27892,g28629);
  and AND2_3385(g28880,g13946,g28639);
  and AND2_3386(g28881,g28612,g9199);
  and AND2_3387(g28892,g14001,g28640);
  and AND2_3388(g28893,g28612,g9245);
  and AND2_3389(g28897,g14016,g28641);
  and AND2_3390(g28898,g28619,g9260);
  and AND2_3391(g28909,g14062,g28642);
  and AND2_3392(g28910,g28612,g9303);
  and AND2_3393(g28914,g14092,g28643);
  and AND2_3394(g28915,g28619,g9323);
  and AND2_3395(g28919,g14107,g28644);
  and AND2_3396(g28923,g28625,g9338);
  and AND2_3397(g28931,g14153,g28645);
  and AND2_3398(g28935,g14177,g28646);
  and AND2_3399(g28936,g28619,g9384);
  and AND2_3400(g28940,g14207,g28647);
  and AND2_3401(g28944,g28625,g9404);
  and AND2_3402(g28948,g14222,g28648);
  and AND2_3403(g28949,g28630,g9419);
  and AND2_3404(g28958,g14268,g28649);
  and AND2_3405(g28962,g14292,g28650);
  and AND2_3406(g28966,g28625,g9481);
  and AND2_3407(g28970,g14322,g28651);
  and AND2_3408(g28971,g28630,g9501);
  and AND2_3409(g28986,g14390,g28652);
  and AND2_3410(g28996,g14414,g28653);
  and AND2_3411(g28997,g28630,g9623);
  and AND2_3412(g29022,g14502,g28655);
  and AND2_3413(g29130,g28397,g22221);
  and AND2_3414(g29174,g29031,g20684);
  and AND2_3415(g29175,g29009,g20687);
  and AND2_3416(g29176,g29097,g20690);
  and AND2_3417(g29180,g28982,g20714);
  and AND2_3418(g29183,g29064,g20739);
  and AND2_3419(g29186,g29063,g20769);
  and AND2_3420(g29188,g29083,g20796);
  and AND2_3421(g29196,g15022,g28741);
  and AND2_3422(g29200,g15096,g28751);
  and AND2_3423(g29203,g15118,g28755);
  and AND2_3424(g29208,g15188,g28764);
  and AND2_3425(g29211,g15210,g28768);
  and AND2_3426(g29217,g15274,g28775);
  and AND2_3427(g29220,g15296,g28779);
  and AND2_3428(g29225,g15366,g28785);
  and AND2_3429(g29229,g9293,g28791);
  and AND2_3430(g29232,g9356,g28796);
  and AND2_3431(g29233,g9374,g28799);
  and AND2_3432(g29234,g9427,g28804);
  and AND2_3433(g29235,g9453,g28807);
  and AND2_3434(g29236,g9471,g28810);
  and AND2_3435(g29238,g9569,g28814);
  and AND2_3436(g29239,g9595,g28817);
  and AND2_3437(g29240,g9613,g28820);
  and AND2_3438(g29241,g9711,g28823);
  and AND2_3439(g29242,g9737,g28826);
  and AND2_3440(g29243,g9857,g28829);
  and AND2_3441(g29248,g28855,g8836);
  and AND2_3442(g29251,g28855,g8856);
  and AND2_3443(g29252,g28859,g8863);
  and AND2_3444(g29255,g28855,g8885);
  and AND2_3445(g29256,g28859,g8894);
  and AND2_3446(g29257,g28863,g8901);
  and AND2_3447(g29259,g28859,g8925);
  and AND2_3448(g29260,g28863,g8934);
  and AND2_3449(g29261,g28867,g8941);
  and AND2_3450(g29262,g28863,g8965);
  and AND2_3451(g29263,g28867,g8974);
  and AND2_3452(g29264,g28867,g8997);
  and AND2_3453(g29284,g29001,g28871);
  and AND2_3454(g29289,g29030,g28883);
  and AND2_3455(g29294,g29053,g28900);
  and AND2_3456(g29300,g29072,g28925);
  and AND2_3457(g29302,g29026,g28928);
  and AND2_3458(g29310,g28978,g28951);
  and AND2_3459(g29312,g29049,g28955);
  and AND2_3460(g29320,g29088,g28972);
  and AND2_3461(g29321,g29008,g28979);
  and AND2_3462(g29323,g29068,g28983);
  and AND2_3463(g29329,g29096,g29002);
  and AND2_3464(g29330,g29038,g29010);
  and AND2_3465(g29332,g29080,g29019);
  and AND2_3466(g29336,g29045,g29023);
  and AND2_3467(g29337,g29103,g29032);
  and AND2_3468(g29338,g29060,g29042);
  and AND2_3469(g29341,g29062,g29046);
  and AND2_3470(g29342,g29107,g29054);
  and AND2_3471(g29344,g29076,g29065);
  and AND2_3472(g29346,g29087,g29077);
  and AND2_3473(g29411,g29090,g21932);
  and AND2_3474(g29464,g29190,g8375);
  and AND2_3475(g29465,g29191,g8424);
  and AND2_3476(g29466,g8587,g29265);
  and AND2_3477(g29467,g29340,g19467);
  and AND2_3478(g29468,g29343,g19490);
  and AND2_3479(g29469,g29345,g19511);
  and AND2_3480(g29470,g29347,g19530);
  and AND2_3481(g29471,g21461,g29266);
  and AND2_3482(g29472,g21461,g29268);
  and AND2_3483(g29473,g21508,g29269);
  and AND2_3484(g29474,g21508,g29271);
  and AND2_3485(g29475,g21544,g29272);
  and AND2_3486(g29476,g21544,g29274);
  and AND2_3487(g29477,g21580,g29275);
  and AND2_3488(g29478,g21580,g29277);
  and AND2_3489(g29479,g21461,g29280);
  and AND2_3490(g29480,g21461,g29282);
  and AND2_3491(g29481,g21508,g29283);
  and AND2_3492(g29482,g21461,g29285);
  and AND2_3493(g29483,g21508,g29286);
  and AND2_3494(g29484,g21544,g29287);
  and AND2_3495(g29485,g21508,g29290);
  and AND2_3496(g29486,g21544,g29291);
  and AND2_3497(g29487,g21580,g29292);
  and AND2_3498(g29488,g21544,g29295);
  and AND2_3499(g29489,g21580,g29296);
  and AND2_3500(g29490,g21580,g29301);
  and AND2_3501(g29502,g29350,g8912);
  and AND2_3502(g29518,g28728,g29360);
  and AND2_3503(g29520,g28731,g29361);
  and AND2_3504(g29521,g28733,g29362);
  and AND2_3505(g29522,g27735,g29363);
  and AND2_3506(g29523,g28737,g29364);
  and AND2_3507(g29524,g28739,g29365);
  and AND2_3508(g29525,g29195,g29366);
  and AND2_3509(g29526,g27741,g29367);
  and AND2_3510(g29527,g28748,g29368);
  and AND2_3511(g29528,g28750,g29369);
  and AND2_3512(g29529,g29199,g29370);
  and AND2_3513(g29531,g29202,g29371);
  and AND2_3514(g29532,g27746,g29372);
  and AND2_3515(g29533,g28762,g29373);
  and AND2_3516(g29534,g29206,g29374);
  and AND2_3517(g29536,g29207,g29375);
  and AND2_3518(g29538,g29210,g29376);
  and AND2_3519(g29539,g27754,g29377);
  and AND2_3520(g29540,g26041,g29378);
  and AND2_3521(g29541,g29214,g29379);
  and AND2_3522(g29543,g29215,g29380);
  and AND2_3523(g29545,g29216,g29381);
  and AND2_3524(g29547,g29219,g29382);
  and AND2_3525(g29548,g28784,g29383);
  and AND2_3526(g29549,g26043,g29384);
  and AND2_3527(g29550,g29222,g29385);
  and AND2_3528(g29553,g29223,g29386);
  and AND2_3529(g29555,g29224,g29387);
  and AND2_3530(g29557,g28789,g29388);
  and AND2_3531(g29558,g28790,g29389);
  and AND2_3532(g29559,g26045,g29390);
  and AND2_3533(g29560,g29227,g29391);
  and AND2_3534(g29562,g29228,g29392);
  and AND2_3535(g29564,g28794,g29393);
  and AND2_3536(g29565,g28795,g29394);
  and AND2_3537(g29566,g26047,g29395);
  and AND2_3538(g29567,g29231,g29396);
  and AND2_3539(g29572,g28802,g29397);
  and AND2_3540(g29573,g28803,g29398);
  and AND2_3541(g29575,g28813,g29402);
  and AND2_3542(g29607,g29193,g11056);
  and AND2_3543(g29610,g29349,g11123);
  and AND2_3544(g29614,g29359,g11182);
  and AND2_3545(g29615,g29245,g11185);
  and AND2_3546(g29619,g29247,g11259);
  and AND2_3547(g29622,g29250,g11327);
  and AND2_3548(g29624,g29254,g11407);
  and AND2_3549(g29625,g29189,g11472);
  and AND2_3550(g29626,g29318,g11478);
  and AND2_3551(g29790,g29491,g10918);
  and AND2_3552(g29792,g29491,g10977);
  and AND2_3553(g29793,g29491,g11063);
  and AND2_3554(g29810,g29748,g22248);
  and AND2_3555(g29811,g29703,g20644);
  and AND2_3556(g29812,g29762,g12223);
  and AND2_3557(g29813,g29760,g13869);
  and AND2_3558(g29814,g29728,g22266);
  and AND2_3559(g29815,g29727,g20662);
  and AND2_3560(g29816,g29759,g13883);
  and AND2_3561(g29817,g29709,g20694);
  and AND2_3562(g29818,g29732,g22293);
  and AND2_3563(g29819,g29751,g22294);
  and AND2_3564(g29820,g29717,g20743);
  and AND2_3565(g29821,g29731,g20746);
  and AND2_3566(g29822,g29705,g22335);
  and AND2_3567(g29827,g29741,g22356);
  and AND2_3568(g29828,g29740,g20802);
  and AND2_3569(g29833,g29725,g20813);
  and AND2_3570(g29834,g29713,g22366);
  and AND2_3571(g29839,g29747,g20827);
  and AND3_256(g29909,g29735,g19420,g19401);
  and AND2_3572(g29910,g29779,g9961);
  and AND2_3573(g29942,g29771,g28877);
  and AND2_3574(g29944,g29782,g28889);
  and AND2_3575(g29945,g29773,g28894);
  and AND2_3576(g29946,g29778,g28906);
  and AND2_3577(g29947,g29785,g28911);
  and AND2_3578(g29948,g29775,g28916);
  and AND2_3579(g29949,g29781,g28932);
  and AND2_3580(g29950,g29788,g28937);
  and AND2_3581(g29951,g29777,g28945);
  and AND2_3582(g29952,g29784,g28959);
  and AND2_3583(g29953,g29791,g28967);
  and AND2_3584(g29954,g29770,g28975);
  and AND2_3585(g29955,g29787,g28993);
  and AND2_3586(g29956,g29780,g28998);
  and AND2_3587(g29957,g29772,g29005);
  and AND2_3588(g29958,g29783,g29027);
  and AND2_3589(g29959,g29774,g29035);
  and AND2_3590(g29960,g29786,g29050);
  and AND2_3591(g29961,g29776,g29057);
  and AND2_3592(g29962,g29789,g29069);
  and AND2_3593(g29963,g29758,g13737);
  and AND2_3594(g29964,g29757,g13786);
  and AND2_3595(g29965,g29756,g11961);
  and AND2_3596(g29966,g29755,g12004);
  and AND2_3597(g29967,g29754,g12066);
  and AND2_3598(g29968,g29765,g12119);
  and AND2_3599(g29969,g29721,g22237);
  and AND2_3600(g29970,g29764,g12178);
  and AND2_3601(g29971,g29763,g13861);
  and AND2_3602(g29980,g29881,g8324);
  and AND2_3603(g29981,g29869,g8330);
  and AND2_3604(g29982,g29893,g8336);
  and AND2_3605(g29983,g29885,g8344);
  and AND2_3606(g29984,g29873,g8351);
  and AND2_3607(g29985,g29897,g8363);
  and AND2_3608(g29986,g29877,g8366);
  and AND2_3609(g29987,g29889,g8369);
  and AND2_3610(g29988,g29881,g8382);
  and AND2_3611(g29989,g29893,g8391);
  and AND2_3612(g29990,g29885,g8397);
  and AND2_3613(g29991,g29901,g8403);
  and AND2_3614(g29992,g12441,g29909);
  and AND2_3615(g29993,g29897,g8411);
  and AND2_3616(g29994,g29889,g8418);
  and AND2_3617(g29995,g29893,g8434);
  and AND2_3618(g29996,g29901,g8443);
  and AND2_3619(g29997,g29918,g22277);
  and AND2_3620(g29998,g29922,g22278);
  and AND2_3621(g29999,g29924,g22279);
  and AND2_3622(g30000,g10767,g29930);
  and AND2_3623(g30001,g29897,g8449);
  and AND2_3624(g30002,g29905,g8455);
  and AND2_3625(g30003,g29901,g8469);
  and AND2_3626(g30004,g29926,g22295);
  and AND2_3627(g30005,g29905,g8478);
  and AND2_3628(g30006,g29928,g22310);
  and AND2_3629(g30007,g29905,g8494);
  and AND2_3630(g30008,g29919,g22334);
  and AND2_3631(g30009,g29929,g22357);
  and AND2_3632(g30077,g29823,g10963);
  and AND2_3633(g30079,g29823,g10988);
  and AND2_3634(g30080,g29829,g10996);
  and AND2_3635(g30081,g29823,g11022);
  and AND2_3636(g30082,g29829,g11036);
  and AND2_3637(g30083,g29835,g11048);
  and AND2_3638(g30085,g29829,g11092);
  and AND2_3639(g30086,g29835,g11108);
  and AND2_3640(g30087,g29840,g11120);
  and AND2_3641(g30088,g29844,g11138);
  and AND2_3642(g30089,g29835,g11160);
  and AND2_3643(g30090,g29840,g11176);
  and AND2_3644(g30091,g29844,g11202);
  and AND2_3645(g30092,g29849,g11205);
  and AND2_3646(g30093,g29853,g11222);
  and AND2_3647(g30094,g29840,g11246);
  and AND2_3648(g30095,g29857,g11265);
  and AND2_3649(g30096,g29844,g11268);
  and AND2_3650(g30097,g29849,g11271);
  and AND2_3651(g30098,g29853,g11284);
  and AND2_3652(g30099,g29861,g11287);
  and AND2_3653(g30100,g29865,g11306);
  and AND2_3654(g30101,g29857,g11341);
  and AND2_3655(g30102,g29849,g11348);
  and AND2_3656(g30103,g29869,g11358);
  and AND2_3657(g30104,g29853,g11361);
  and AND2_3658(g30105,g29861,g11364);
  and AND2_3659(g30106,g29865,g11379);
  and AND2_3660(g30107,g29873,g11382);
  and AND2_3661(g30108,g29877,g11401);
  and AND2_3662(g30109,g29857,g11411);
  and AND2_3663(g30110,g29881,g11417);
  and AND2_3664(g30111,g29869,g11425);
  and AND2_3665(g30112,g29861,g11432);
  and AND2_3666(g30113,g29885,g11444);
  and AND2_3667(g30114,g29865,g11447);
  and AND2_3668(g30115,g29873,g11450);
  and AND2_3669(g30116,g29921,g22236);
  and AND2_3670(g30117,g29877,g11465);
  and AND2_3671(g30118,g29889,g11468);
  and AND2_3672(g30123,g30070,g20641);
  and AND2_3673(g30127,g30065,g20719);
  and AND2_3674(g30128,g30062,g20722);
  and AND2_3675(g30129,g30071,g20725);
  and AND2_3676(g30131,g30059,g20749);
  and AND2_3677(g30132,g30068,g20776);
  and AND2_3678(g30133,g30067,g20799);
  and AND2_3679(g30138,g30069,g20816);
  and AND2_3680(g30216,g30036,g8921);
  and AND2_3681(g30217,g30036,g8955);
  and AND2_3682(g30218,g30040,g8961);
  and AND2_3683(g30219,g30036,g8980);
  and AND2_3684(g30220,g30040,g8987);
  and AND2_3685(g30221,g30044,g8993);
  and AND2_3686(g30222,g30040,g9010);
  and AND2_3687(g30223,g30044,g9016);
  and AND2_3688(g30224,g30048,g9022);
  and AND2_3689(g30225,g30044,g9035);
  and AND2_3690(g30226,g30048,g9041);
  and AND2_3691(g30227,g30048,g9058);
  and AND2_3692(g30327,g30187,g8321);
  and AND2_3693(g30330,g30195,g8333);
  and AND2_3694(g30333,g30191,g8341);
  and AND2_3695(g30334,g30203,g8347);
  and AND2_3696(g30337,g30199,g8354);
  and AND2_3697(g30340,g30207,g8372);
  and AND2_3698(g30345,g30195,g8388);
  and AND2_3699(g30348,g30203,g8400);
  and AND2_3700(g30351,g30199,g8408);
  and AND2_3701(g30352,g30211,g8414);
  and AND2_3702(g30355,g30207,g8421);
  and AND2_3703(g30361,g30203,g8440);
  and AND2_3704(g30364,g30211,g8452);
  and AND2_3705(g30367,g30207,g8460);
  and AND2_3706(g30372,g8594,g30228);
  and AND2_3707(g30374,g30211,g8475);
  and AND2_3708(g30387,g30229,g8888);
  and AND2_3709(g30388,g30229,g8918);
  and AND2_3710(g30389,g30233,g8928);
  and AND2_3711(g30390,g30229,g8952);
  and AND2_3712(g30391,g30233,g8958);
  and AND2_3713(g30392,g30237,g8968);
  and AND2_3714(g30393,g30233,g8984);
  and AND2_3715(g30394,g30237,g8990);
  and AND2_3716(g30395,g30241,g9000);
  and AND2_3717(g30396,g30237,g9013);
  and AND2_3718(g30397,g30241,g9019);
  and AND2_3719(g30398,g30241,g9038);
  and AND2_3720(g30407,g30134,g10991);
  and AND2_3721(g30409,g30134,g11025);
  and AND2_3722(g30410,g30139,g11028);
  and AND2_3723(g30411,g30143,g11039);
  and AND2_3724(g30436,g30134,g11079);
  and AND2_3725(g30437,g30139,g11082);
  and AND2_3726(g30438,g30147,g11085);
  and AND2_3727(g30440,g30143,g11095);
  and AND2_3728(g30441,g30151,g11098);
  and AND2_3729(g30442,g30155,g11111);
  and AND2_3730(g30444,g30139,g11132);
  and AND2_3731(g30445,g30147,g11135);
  and AND2_3732(g30447,g30143,g11145);
  and AND2_3733(g30448,g30151,g11148);
  and AND2_3734(g30449,g30159,g11151);
  and AND2_3735(g30451,g30155,g11163);
  and AND2_3736(g30452,g30163,g11166);
  and AND2_3737(g30453,g30167,g11179);
  and AND2_3738(g30454,g30147,g11199);
  and AND2_3739(g30457,g30151,g11216);
  and AND2_3740(g30458,g30159,g11219);
  and AND2_3741(g30460,g30155,g11231);
  and AND2_3742(g30461,g30163,g11234);
  and AND2_3743(g30462,g30171,g11237);
  and AND2_3744(g30464,g30167,g11249);
  and AND2_3745(g30465,g30175,g11252);
  and AND2_3746(g30467,g30179,g11274);
  and AND2_3747(g30469,g30159,g11281);
  and AND2_3748(g30472,g30163,g11300);
  and AND2_3749(g30473,g30171,g11303);
  and AND2_3750(g30475,g30167,g11315);
  and AND2_3751(g30476,g30175,g11318);
  and AND2_3752(g30477,g30183,g11321);
  and AND2_3753(g30478,g30187,g11344);
  and AND2_3754(g30481,g30179,g11351);
  and AND2_3755(g30484,g30191,g11367);
  and AND2_3756(g30486,g30171,g11376);
  and AND2_3757(g30489,g30175,g11395);
  and AND2_3758(g30490,g30183,g11398);
  and AND2_3759(g30492,g30187,g11414);
  and AND2_3760(g30495,g30179,g11422);
  and AND2_3761(g30496,g30195,g11428);
  and AND2_3762(g30499,g30191,g11435);
  and AND2_3763(g30502,g30199,g11453);
  and AND2_3764(g30504,g30183,g11462);
  and AND2_3765(g30696,g30383,g10943);
  and AND2_3766(g30697,g30383,g11011);
  and AND2_3767(g30698,g30383,g11126);
  and AND2_3768(g30728,g30605,g22252);
  and AND2_3769(g30735,g30629,g22268);
  and AND2_3770(g30736,g30584,g20669);
  and AND2_3771(g30743,g30610,g22283);
  and AND2_3772(g30744,g30609,g20697);
  and AND2_3773(g30750,g30593,g20729);
  and AND2_3774(g30754,g30614,g22313);
  and AND2_3775(g30755,g30632,g22314);
  and AND2_3776(g30757,g30601,g20780);
  and AND2_3777(g30758,g30613,g20783);
  and AND2_3778(g30759,g30588,g22360);
  and AND2_3779(g30760,g30622,g22379);
  and AND2_3780(g30761,g30621,g20822);
  and AND2_3781(g30762,g30608,g20830);
  and AND2_3782(g30763,g30597,g22386);
  and AND2_3783(g30764,g30628,g20837);
  and AND3_257(g30766,g30617,g19457,g19431);
  and AND2_3784(g30916,g30785,g22251);
  and AND2_3785(g30917,g12446,g30766);
  and AND2_3786(g30918,g30780,g22296);
  and AND2_3787(g30919,g30786,g22297);
  and AND2_3788(g30920,g30787,g22298);
  and AND2_3789(g30921,g10773,g30791);
  and AND2_3790(g30922,g30788,g22315);
  and AND2_3791(g30923,g30789,g22338);
  and AND2_3792(g30924,g30783,g22359);
  and AND2_3793(g30925,g30790,g22380);
  and AND2_3794(g30944,g30935,g20666);
  and AND2_3795(g30945,g30931,g20754);
  and AND2_3796(g30946,g30930,g20757);
  and AND2_3797(g30947,g30936,g20760);
  and AND2_3798(g30948,g30929,g20786);
  and AND2_3799(g30949,g30933,g20806);
  and AND2_3800(g30950,g30932,g20819);
  and AND2_3801(g30951,g30934,g20833);
  and AND2_3802(g30953,g8605,g30952);
  or OR2_0(g9144,g2986,g5389);
  or OR2_1(g10778,g2929,g8022);
  or OR2_2(g12377,g7553,g11059);
  or OR2_3(g12407,g7573,g10779);
  or OR2_4(g12886,g9534,g3398);
  or OR2_5(g12926,g9676,g3554);
  or OR2_6(g12955,g9822,g3710);
  or OR2_7(g12984,g9968,g3866);
  or OR2_8(g16539,g15880,g14657);
  or OR2_9(g16571,g15913,g14691);
  or OR2_10(g16595,g15942,g14725);
  or OR2_11(g16615,g15971,g14753);
  or OR2_12(g17973,g11623,g15659);
  or OR2_13(g19181,g17729,g17979);
  or OR2_14(g19186,g18419,g17887);
  or OR2_15(g19187,g18419,g17729);
  or OR2_16(g19188,g17830,g18096);
  or OR2_17(g19191,g17807,g17887);
  or OR2_18(g19192,g18183,g18270);
  or OR2_19(g19193,g18492,g17998);
  or OR2_20(g19194,g18492,g17830);
  or OR2_21(g19195,g17942,g18212);
  or OR2_22(g19200,g18346,g18424);
  or OR2_23(g19201,g18183,g18424);
  or OR2_24(g19202,g17919,g17998);
  or OR2_25(g19203,g18290,g18363);
  or OR2_26(g19204,g18556,g18115);
  or OR2_27(g19205,g18556,g17942);
  or OR2_28(g19206,g18053,g18319);
  or OR2_29(g19209,g18079,g18346);
  or OR2_30(g19210,g18079,g18183);
  or OR2_31(g19211,g18441,g18497);
  or OR2_32(g19212,g18290,g18497);
  or OR2_33(g19213,g18030,g18115);
  or OR2_34(g19214,g18383,g18458);
  or OR2_35(g19215,g18606,g18231);
  or OR2_36(g19216,g18606,g18053);
  or OR2_37(g19221,g18270,g18346);
  or OR2_38(g19222,g18195,g18441);
  or OR2_39(g19223,g18195,g18290);
  or OR2_40(g19224,g18514,g18561);
  or OR2_41(g19225,g18383,g18561);
  or OR2_42(g19226,g18147,g18231);
  or OR2_43(g19227,g18478,g18531);
  or OR3_0(II25477,g17024,g17000,g16992);
  or OR3_1(g19230,g16985,g16965,II25477);
  or OR2_44(g19231,g18363,g18441);
  or OR2_45(g19232,g18302,g18514);
  or OR2_46(g19233,g18302,g18383);
  or OR2_47(g19234,g18578,g18611);
  or OR2_48(g19235,g18478,g18611);
  or OR3_2(II25495,g17158,g17137,g17115);
  or OR3_3(g19240,g17083,g17050,II25495);
  or OR2_49(g19242,g14244,g16501);
  or OR3_4(II25500,g17058,g17030,g17016);
  or OR3_5(g19243,g16995,g16986,II25500);
  or OR2_50(g19244,g18458,g18514);
  or OR2_51(g19245,g18395,g18578);
  or OR2_52(g19246,g18395,g18478);
  or OR2_53(g19250,g17729,g17807);
  or OR3_6(II25516,g17173,g17160,g17142);
  or OR3_7(g19253,g17121,g17085,II25516);
  or OR2_54(g19255,g14366,g16523);
  or OR3_8(II25521,g17093,g17064,g17046);
  or OR3_9(g19256,g17019,g16996,II25521);
  or OR2_55(g19257,g18531,g18578);
  or OR2_56(g19263,g17887,g17979);
  or OR2_57(g19264,g17830,g17919);
  or OR3_10(II25549,g17190,g17175,g17165);
  or OR3_11(g19266,g17148,g17123,II25549);
  or OR2_58(g19268,g14478,g16554);
  or OR3_12(II25554,g17131,g17099,g17080);
  or OR3_13(g19269,g17049,g17020,II25554);
  or OR3_14(g19275,g16867,g16515,g19001);
  or OR2_59(g19278,g17998,g18096);
  or OR2_60(g19279,g17942,g18030);
  or OR3_15(II25588,g17201,g17192,g17180);
  or OR3_16(g19281,g17171,g17150,II25588);
  or OR2_61(g19283,g14565,g16586);
  or OR3_17(g19294,g16895,g16546,g16507);
  or OR2_62(g19297,g18115,g18212);
  or OR2_63(g19298,g18053,g18147);
  or OR3_18(g19312,g16924,g16578,g16529);
  or OR2_64(g19315,g18231,g18319);
  or OR3_19(g19333,g16954,g16602,g16560);
  or OR2_65(g19450,g14837,g16682);
  or OR2_66(g19477,g14910,g16708);
  or OR2_67(g19500,g14991,g16739);
  or OR3_20(g19503,g16884,g16697,g16665);
  or OR2_68(g19521,g15080,g16781);
  or OR3_21(g19522,g16913,g16728,g16686);
  or OR3_22(g19532,g16943,g16770,g16712);
  or OR3_23(g19542,g16974,g16797,g16743);
  or OR3_24(II26429,g17979,g17887,g17807);
  or OR3_25(g19981,g17729,g18419,II26429);
  or OR3_26(II26455,g18424,g18346,g18270);
  or OR3_27(g20015,g18183,g18079,II26455);
  or OR3_28(II26461,g18096,g17998,g17919);
  or OR3_29(g20019,g17830,g18492,II26461);
  or OR3_30(II26491,g18497,g18441,g18363);
  or OR3_31(g20057,g18290,g18195,II26491);
  or OR3_32(II26497,g18212,g18115,g18030);
  or OR3_33(g20061,g17942,g18556,II26497);
  or OR3_34(II26532,g18561,g18514,g18458);
  or OR3_35(g20098,g18383,g18302,II26532);
  or OR3_36(II26538,g18319,g18231,g18147);
  or OR3_37(g20102,g18053,g18606,II26538);
  or OR3_38(II26571,g18611,g18578,g18531);
  or OR3_39(g20123,g18478,g18395,II26571);
  or OR3_40(g21120,g19484,g16515,g14071);
  or OR3_41(g21139,g19505,g16546,g14186);
  or OR3_42(g21159,g19524,g16578,g14301);
  or OR3_43(g21179,g19534,g16602,g14423);
  or OR3_44(g21244,g19578,g16697,g14776);
  or OR3_45(g21253,g19608,g16728,g14811);
  or OR3_46(g21261,g19641,g16770,g14863);
  or OR3_47(g21269,g19681,g16797,g14936);
  or OR3_48(g21501,g20522,g16867,g14071);
  or OR3_49(g21536,g20522,g19484,g19001);
  or OR3_50(g21540,g20542,g16895,g14186);
  or OR3_51(g21572,g20542,g19505,g16507);
  or OR3_52(g21576,g19067,g16924,g14301);
  or OR3_53(g21605,g19067,g19524,g16529);
  or OR3_54(g21609,g19084,g16954,g14423);
  or OR3_55(g21634,g19084,g19534,g16560);
  or OR3_56(g21774,g19121,g16884,g14776);
  or OR3_57(g21787,g19121,g19578,g16665);
  or OR3_58(II28305,g20197,g20177,g20145);
  or OR3_59(g21788,g20117,g20094,II28305);
  or OR3_60(g21789,g19128,g16913,g14811);
  or OR3_61(II28318,g19092,g19088,g19079);
  or OR4_0(g21799,g16505,g20538,g18994,II28318);
  or OR4_1(g21800,g18665,g20270,g20248,g18647);
  or OR3_62(g21801,g19128,g19608,g16686);
  or OR3_63(II28323,g20227,g20211,g20183);
  or OR3_64(g21802,g20147,g20119,II28323);
  or OR3_65(g21803,g19135,g16943,g14863);
  or OR4_2(g21806,g20116,g20093,g18547,g19097);
  or OR3_66(II28330,g19099,g19094,g19089);
  or OR4_3(g21807,g16527,g19063,g19007,II28330);
  or OR4_4(g21808,g18688,g20282,g20271,g18650);
  or OR3_67(g21809,g19135,g19641,g16712);
  or OR3_68(II28335,g20254,g20241,g20217);
  or OR3_69(g21810,g20185,g20149,II28335);
  or OR3_70(g21811,g19138,g16974,g14936);
  or OR4_5(g21813,g20146,g20118,g18597,g19104);
  or OR3_71(II28341,g19106,g19101,g19095);
  or OR4_6(g21814,g16558,g19080,g16513,II28341);
  or OR4_7(g21815,g18717,g20293,g20283,g18654);
  or OR3_72(g21816,g19138,g19681,g16743);
  or OR3_73(II28346,g20277,g20268,g20247);
  or OR3_74(g21817,g20219,g20187,II28346);
  or OR4_8(g21819,g20184,g20148,g18629,g19109);
  or OR3_75(II28351,g19111,g19108,g19102);
  or OR4_9(g21820,g16590,g19090,g16535,II28351);
  or OR4_10(g21821,g18753,g20309,g20294,g18668);
  or OR4_11(g21823,g20218,g20186,g18638,g19116);
  or OR3_76(II28365,g20280,g18652,g18649);
  or OR3_77(g21844,g20222,g18645,II28365);
  or OR3_78(II28369,g20291,g18666,g18653);
  or OR3_79(g21846,g20249,g18648,II28369);
  or OR3_80(II28374,g20307,g18689,g18667);
  or OR3_81(g21849,g20272,g18651,II28374);
  or OR3_82(II28380,g20326,g18718,g18690);
  or OR3_83(g21856,g20284,g18655,II28380);
  or OR2_69(g22175,g16075,g20842);
  or OR2_70(g22190,g16113,g20850);
  or OR2_71(g22199,g16164,g20858);
  or OR2_72(g22205,g16223,g20866);
  or OR4_12(g22811,g562,g559,g12451,g21851);
  or OR3_84(g23052,g21800,g21788,g21844);
  or OR3_85(g23071,g21808,g21802,g21846);
  or OR3_86(g23084,g21815,g21810,g21849);
  or OR2_73(g23089,g21806,g21799);
  or OR3_87(g23100,g21821,g21817,g21856);
  or OR2_74(g23107,g21813,g21807);
  or OR2_75(g23120,g21819,g21814);
  or OR2_76(g23129,g21823,g21820);
  or OR2_77(g23319,g14493,g22385);
  or OR2_78(g23688,g23106,g21906);
  or OR2_79(g23742,g23119,g21920);
  or OR2_80(g23797,g23128,g21938);
  or OR2_81(g23850,g23139,g20647);
  or OR2_82(g23919,g22666,g23140);
  or OR2_83(g24239,g19387,g22401);
  or OR2_84(g24244,g14144,g22317);
  or OR2_85(g24245,g19417,g22402);
  or OR2_86(g24252,g14259,g22342);
  or OR2_87(g24254,g19454,g22403);
  or OR2_88(g24257,g14381,g22365);
  or OR2_89(g24258,g19481,g22404);
  or OR2_90(g24633,g24094,g20842);
  or OR2_91(g24653,g24095,g20850);
  or OR2_92(g24672,g24097,g20858);
  or OR2_93(g24691,g24103,g20866);
  or OR2_94(g24890,g23639,g23144);
  or OR2_95(g24909,g23726,g23142);
  or OR2_96(g24925,g23772,g23141);
  or OR2_97(g24965,g23922,g23945);
  or OR2_98(g24978,g23954,g23974);
  or OR2_99(g24989,g23983,g24004);
  or OR2_100(g25000,g24013,g24038);
  or OR2_101(g25183,g24958,g24893);
  or OR2_102(g25186,g24969,g24916);
  or OR2_103(g25190,g24982,g24933);
  or OR2_104(g25195,g24993,g24945);
  or OR2_105(g25489,g24795,g16466);
  or OR2_106(g25490,g24759,g23146);
  or OR2_107(g25520,g24813,g23145);
  or OR2_108(g25566,g24843,g23143);
  or OR2_109(g26320,g25852,g25870);
  or OR2_110(g26367,g25873,g25882);
  or OR2_111(g26410,g25885,g25887);
  or OR2_112(g26451,g25890,g25892);
  or OR2_113(g26974,g26157,g23147);
  or OR3_88(g27113,g1248,g1245,g26534);
  or OR2_114(g28501,g27738,g25764);
  or OR2_115(g28512,g26481,g27738);
  or OR2_116(g28529,g27743,g25818);
  or OR2_117(g28540,g26497,g27743);
  or OR2_118(g28556,g27751,g25853);
  or OR2_119(g28567,g26512,g27751);
  or OR2_120(g28584,g27756,g25874);
  or OR2_121(g28595,g26520,g27756);
  or OR3_89(g29348,g1942,g1939,g29113);
  or OR3_90(g30305,g2636,g2633,g30072);
  nand NAND2_0(II15167,g2981,g2874);
  nand NAND2_1(II15168,g2981,II15167);
  nand NAND2_2(II15169,g2874,II15167);
  nand NAND2_3(g7855,II15168,II15169);
  nand NAND2_4(II15183,g2975,g2978);
  nand NAND2_5(II15184,g2975,II15183);
  nand NAND2_6(II15185,g2978,II15183);
  nand NAND2_7(g7875,II15184,II15185);
  nand NAND2_8(II15190,g2956,g2959);
  nand NAND2_9(II15191,g2956,II15190);
  nand NAND2_10(II15192,g2959,II15190);
  nand NAND2_11(g7876,II15191,II15192);
  nand NAND2_12(II15204,g2969,g2972);
  nand NAND2_13(II15205,g2969,II15204);
  nand NAND2_14(II15206,g2972,II15204);
  nand NAND2_15(g7895,II15205,II15206);
  nand NAND2_16(II15211,g2947,g2953);
  nand NAND2_17(II15212,g2947,II15211);
  nand NAND2_18(II15213,g2953,II15211);
  nand NAND2_19(g7896,II15212,II15213);
  nand NAND2_20(II15237,g2963,g2966);
  nand NAND2_21(II15238,g2963,II15237);
  nand NAND2_22(II15239,g2966,II15237);
  nand NAND2_23(g7922,II15238,II15239);
  nand NAND2_24(II15244,g2941,g2944);
  nand NAND2_25(II15245,g2941,II15244);
  nand NAND2_26(II15246,g2944,II15244);
  nand NAND2_27(g7923,II15245,II15246);
  nand NAND2_28(II15276,g2935,g2938);
  nand NAND2_29(II15277,g2935,II15276);
  nand NAND2_30(II15278,g2938,II15276);
  nand NAND2_31(g7970,II15277,II15278);
  nand NAND4_0(g8381,g8182,g8120,g8044,g7989);
  nand NAND2_32(g8533,g3398,g3366);
  nand NAND2_33(g8547,g3398,g3366);
  nand NAND2_34(g8550,g3554,g3522);
  nand NAND2_35(g8560,g3554,g3522);
  nand NAND2_36(g8563,g3710,g3678);
  nand NAND2_37(g8571,g3710,g3678);
  nand NAND2_38(g8574,g3866,g3834);
  nand NAND2_39(g8577,g3866,g3834);
  nand NAND2_40(II16879,g4203,g3998);
  nand NAND2_41(II16880,g4203,II16879);
  nand NAND2_42(II16881,g3998,II16879);
  nand NAND2_43(g9883,II16880,II16881);
  nand NAND2_44(II16965,g4734,g4452);
  nand NAND2_45(II16966,g4734,II16965);
  nand NAND2_46(II16967,g4452,II16965);
  nand NAND2_47(g10003,II16966,II16967);
  nand NAND2_48(g10038,g7772,g3366);
  nand NAND2_49(II17059,g6637,g6309);
  nand NAND2_50(II17060,g6637,II17059);
  nand NAND2_51(II17061,g6309,II17059);
  nand NAND2_52(g10095,II17060,II17061);
  nand NAND2_53(g10147,g7788,g3522);
  nand NAND2_54(II17149,g7465,g7142);
  nand NAND2_55(II17150,g7465,II17149);
  nand NAND2_56(II17151,g7142,II17149);
  nand NAND2_57(g10185,II17150,II17151);
  nand NAND2_58(g10252,g7802,g3678);
  nand NAND2_59(g10354,g7815,g3834);
  nand NAND2_60(g10649,g3398,g6912);
  nand NAND2_61(g10676,g3398,g6678);
  nand NAND2_62(g10677,g3398,g6912);
  nand NAND2_63(g10679,g3554,g7162);
  nand NAND2_64(g10703,g3398,g6678);
  nand NAND2_65(g10705,g3554,g6980);
  nand NAND2_66(g10706,g3554,g7162);
  nand NAND2_67(g10708,g3710,g7358);
  nand NAND2_68(g10723,g3554,g6980);
  nand NAND2_69(g10725,g3710,g7230);
  nand NAND2_70(g10726,g3710,g7358);
  nand NAND2_71(g10728,g3866,g7488);
  nand NAND2_72(g10744,g3710,g7230);
  nand NAND2_73(g10746,g3866,g7426);
  nand NAND2_74(g10747,g3866,g7488);
  nand NAND2_75(g10763,g3866,g7426);
  nand NAND2_76(II18106,g7875,g7855);
  nand NAND2_77(II18107,g7875,II18106);
  nand NAND2_78(II18108,g7855,II18106);
  nand NAND2_79(g11188,II18107,II18108);
  nand NAND2_80(II18113,g3997,g8181);
  nand NAND2_81(II18114,g3997,II18113);
  nand NAND2_82(II18115,g8181,II18113);
  nand NAND2_83(g11189,II18114,II18115);
  nand NAND2_84(II18190,g7922,g7895);
  nand NAND2_85(II18191,g7922,II18190);
  nand NAND2_86(II18192,g7895,II18190);
  nand NAND2_87(g11262,II18191,II18192);
  nand NAND2_88(II18197,g7896,g7876);
  nand NAND2_89(II18198,g7896,II18197);
  nand NAND2_90(II18199,g7876,II18197);
  nand NAND2_91(g11263,II18198,II18199);
  nand NAND2_92(II18204,g7975,g4202);
  nand NAND2_93(II18205,g7975,II18204);
  nand NAND2_94(II18206,g4202,II18204);
  nand NAND2_95(g11264,II18205,II18206);
  nand NAND2_96(II18280,g7970,g7923);
  nand NAND2_97(II18281,g7970,II18280);
  nand NAND2_98(II18282,g7923,II18280);
  nand NAND2_99(g11330,II18281,II18282);
  nand NAND2_100(II18287,g8256,g8102);
  nand NAND2_101(II18288,g8256,II18287);
  nand NAND2_102(II18289,g8102,II18287);
  nand NAND2_103(g11331,II18288,II18289);
  nand NAND2_104(II18368,g4325,g4093);
  nand NAND2_105(II18369,g4325,II18368);
  nand NAND2_106(II18370,g4093,II18368);
  nand NAND2_107(g11410,II18369,II18370);
  nand NAND2_108(g11617,g8313,g2883);
  nand NAND2_109(II18799,g11410,g11331);
  nand NAND2_110(II18800,g11410,II18799);
  nand NAND2_111(II18801,g11331,II18799);
  nand NAND2_112(g11621,II18800,II18801);
  nand NAND2_113(g11661,g9534,g3366);
  nand NAND2_114(g11662,g9534,g3366);
  nand NAND2_115(g11672,g9534,g3366);
  nand NAND2_116(g11673,g9676,g3522);
  nand NAND2_117(g11674,g9676,g3522);
  nand NAND2_118(g11683,g9534,g3366);
  nand NAND2_119(g11684,g9676,g3522);
  nand NAND2_120(g11685,g9822,g3678);
  nand NAND2_121(g11686,g9822,g3678);
  nand NAND2_122(g11691,g9534,g3366);
  nand NAND2_123(g11692,g9676,g3522);
  nand NAND2_124(g11693,g9822,g3678);
  nand NAND2_125(g11694,g9968,g3834);
  nand NAND2_126(g11695,g9968,g3834);
  nand NAND2_127(g11696,g9534,g3366);
  nand NAND2_128(g11698,g9676,g3522);
  nand NAND2_129(g11699,g9822,g3678);
  nand NAND2_130(g11700,g9968,g3834);
  nand NAND2_131(g11701,g9534,g3366);
  nand NAND2_132(g11702,g9676,g3522);
  nand NAND2_133(g11704,g9822,g3678);
  nand NAND2_134(g11705,g9968,g3834);
  nand NAND2_135(g11707,g9534,g3366);
  nand NAND2_136(g11708,g9534,g3366);
  nand NAND2_137(g11709,g9676,g3522);
  nand NAND2_138(g11710,g9822,g3678);
  nand NAND2_139(g11712,g9968,g3834);
  nand NAND2_140(g11713,g10481,g9144);
  nand NAND2_141(g11716,g9534,g3366);
  nand NAND2_142(g11717,g9676,g3522);
  nand NAND2_143(g11718,g9676,g3522);
  nand NAND2_144(g11719,g9822,g3678);
  nand NAND2_145(g11720,g9968,g3834);
  nand NAND2_146(g11721,g9534,g3366);
  nand NAND2_147(g11722,g9676,g3522);
  nand NAND2_148(g11723,g9822,g3678);
  nand NAND2_149(g11724,g9822,g3678);
  nand NAND2_150(g11725,g9968,g3834);
  nand NAND2_151(g11726,g9676,g3522);
  nand NAND2_152(g11727,g9822,g3678);
  nand NAND2_153(g11728,g9968,g3834);
  nand NAND2_154(g11729,g9968,g3834);
  nand NAND2_155(g11730,g9822,g3678);
  nand NAND2_156(g11731,g9968,g3834);
  nand NAND2_157(g11733,g9968,g3834);
  nand NAND2_158(g12433,g2879,g10778);
  nand NAND2_159(g12486,g8278,g6448);
  nand NAND2_160(g12503,g8278,g5438);
  nand NAND2_161(g12506,g8287,g6713);
  nand NAND2_162(g12520,g8287,g5473);
  nand NAND2_163(g12523,g8296,g7015);
  nand NAND2_164(g12535,g8296,g5512);
  nand NAND2_165(g12538,g8305,g7265);
  nand NAND2_166(g12544,g8305,g5556);
  nand NAND2_167(II20031,g10003,g9883);
  nand NAND2_168(II20032,g10003,II20031);
  nand NAND2_169(II20033,g9883,II20031);
  nand NAND2_170(g12988,II20032,II20033);
  nand NAND2_171(II20048,g10185,g10095);
  nand NAND2_172(II20049,g10185,II20048);
  nand NAND2_173(II20050,g10095,II20048);
  nand NAND2_174(g12999,II20049,II20050);
  nand NAND2_175(g13020,g9534,g6912);
  nand NAND2_176(g13021,g9534,g6912);
  nand NAND2_177(g13026,g9534,g6678);
  nand NAND2_178(g13027,g9534,g6912);
  nand NAND2_179(g13028,g9534,g6678);
  nand NAND2_180(g13029,g9676,g7162);
  nand NAND2_181(g13030,g9676,g7162);
  nand NAND2_182(g13034,g9534,g6678);
  nand NAND2_183(g13035,g9534,g6912);
  nand NAND2_184(g13037,g9676,g6980);
  nand NAND2_185(g13038,g9676,g7162);
  nand NAND2_186(g13039,g9676,g6980);
  nand NAND2_187(g13040,g9822,g7358);
  nand NAND2_188(g13041,g9822,g7358);
  nand NAND2_189(g13044,g9534,g6678);
  nand NAND2_190(g13045,g9534,g6912);
  nand NAND2_191(g13047,g9676,g6980);
  nand NAND2_192(g13048,g9676,g7162);
  nand NAND2_193(g13050,g9822,g7230);
  nand NAND2_194(g13051,g9822,g7358);
  nand NAND2_195(g13052,g9822,g7230);
  nand NAND2_196(g13053,g9968,g7488);
  nand NAND2_197(g13054,g9968,g7488);
  nand NAND2_198(g13058,g9534,g6678);
  nand NAND2_199(g13059,g9534,g6912);
  nand NAND2_200(g13061,g9676,g6980);
  nand NAND2_201(g13062,g9676,g7162);
  nand NAND2_202(g13064,g9822,g7230);
  nand NAND2_203(g13065,g9822,g7358);
  nand NAND2_204(g13067,g9968,g7426);
  nand NAND2_205(g13068,g9968,g7488);
  nand NAND2_206(g13069,g9968,g7426);
  nand NAND2_207(g13071,g9534,g6678);
  nand NAND2_208(g13072,g9534,g6912);
  nand NAND2_209(g13074,g9676,g6980);
  nand NAND2_210(g13075,g9676,g7162);
  nand NAND2_211(g13077,g9822,g7230);
  nand NAND2_212(g13078,g9822,g7358);
  nand NAND2_213(g13080,g9968,g7426);
  nand NAND2_214(g13081,g9968,g7488);
  nand NAND2_215(g13087,g9534,g6678);
  nand NAND2_216(g13088,g9534,g6912);
  nand NAND2_217(g13089,g9534,g6912);
  nand NAND2_218(g13090,g9676,g6980);
  nand NAND2_219(g13091,g9676,g7162);
  nand NAND2_220(g13093,g9822,g7230);
  nand NAND2_221(g13094,g9822,g7358);
  nand NAND2_222(g13096,g9968,g7426);
  nand NAND2_223(g13097,g9968,g7488);
  nand NAND2_224(g13098,g9534,g6678);
  nand NAND2_225(g13099,g9534,g6912);
  nand NAND2_226(g13100,g9534,g6678);
  nand NAND2_227(g13102,g9676,g6980);
  nand NAND2_228(g13103,g9676,g7162);
  nand NAND2_229(g13104,g9676,g7162);
  nand NAND2_230(g13105,g9822,g7230);
  nand NAND2_231(g13106,g9822,g7358);
  nand NAND2_232(g13108,g9968,g7426);
  nand NAND2_233(g13109,g9968,g7488);
  nand NAND2_234(g13112,g9534,g6678);
  nand NAND2_235(g13113,g9534,g6912);
  nand NAND2_236(g13114,g9676,g6980);
  nand NAND2_237(g13115,g9676,g7162);
  nand NAND2_238(g13116,g9676,g6980);
  nand NAND2_239(g13118,g9822,g7230);
  nand NAND2_240(g13119,g9822,g7358);
  nand NAND2_241(g13120,g9822,g7358);
  nand NAND2_242(g13121,g9968,g7426);
  nand NAND2_243(g13122,g9968,g7488);
  nand NAND2_244(g13123,g9534,g6678);
  nand NAND2_245(g13125,g9676,g6980);
  nand NAND2_246(g13126,g9676,g7162);
  nand NAND2_247(g13127,g9822,g7230);
  nand NAND2_248(g13128,g9822,g7358);
  nand NAND2_249(g13129,g9822,g7230);
  nand NAND2_250(g13131,g9968,g7426);
  nand NAND2_251(g13132,g9968,g7488);
  nand NAND2_252(g13133,g9968,g7488);
  nand NAND2_253(g13134,g9676,g6980);
  nand NAND2_254(g13136,g9822,g7230);
  nand NAND2_255(g13137,g9822,g7358);
  nand NAND2_256(g13138,g9968,g7426);
  nand NAND2_257(g13139,g9968,g7488);
  nand NAND2_258(g13140,g9968,g7426);
  nand NAND2_259(g13142,g9822,g7230);
  nand NAND2_260(g13144,g9968,g7426);
  nand NAND2_261(g13145,g9968,g7488);
  nand NAND2_262(g13146,g9968,g7426);
  nand NAND2_263(g13147,g8278,g3306);
  nand NAND2_264(g13150,g8287,g3462);
  nand NAND2_265(g13156,g8296,g3618);
  nand NAND2_266(g13165,g8305,g3774);
  nand NAND2_267(g13245,g10779,g7901);
  nand NAND2_268(g13305,g8317,g2993);
  nand NAND2_269(II20429,g11262,g11188);
  nand NAND2_270(II20430,g11262,II20429);
  nand NAND2_271(II20431,g11188,II20429);
  nand NAND2_272(g13348,II20430,II20431);
  nand NAND2_273(II20465,g11330,g11263);
  nand NAND2_274(II20466,g11330,II20465);
  nand NAND2_275(II20467,g11263,II20465);
  nand NAND2_276(g13370,II20466,II20467);
  nand NAND2_277(II20504,g11264,g11189);
  nand NAND2_278(II20505,g11264,II20504);
  nand NAND2_279(II20506,g11189,II20504);
  nand NAND2_280(g13399,II20505,II20506);
  nand NAND2_281(g13476,g12565,g3254);
  nand NAND2_282(g13478,g12611,g3410);
  nand NAND2_283(g13482,g12657,g3566);
  nand NAND2_284(g13494,g12565,g3254);
  nand NAND2_285(g13495,g12611,g3410);
  nand NAND2_286(g13497,g12657,g3566);
  nand NAND2_287(g13501,g12711,g3722);
  nand NAND2_288(II20743,g11621,g13399);
  nand NAND2_289(II20744,g11621,II20743);
  nand NAND2_290(II20745,g13399,II20743);
  nand NAND2_291(g13507,II20744,II20745);
  nand NAND2_292(g13510,g12565,g3254);
  nand NAND2_293(g13511,g12611,g3410);
  nand NAND2_294(g13512,g12657,g3566);
  nand NAND2_295(g13514,g12711,g3722);
  nand NAND2_296(g13518,g12565,g3254);
  nand NAND2_297(g13524,g12611,g3410);
  nand NAND2_298(g13525,g12657,g3566);
  nand NAND2_299(g13526,g12711,g3722);
  nand NAND2_300(g13528,g12565,g3254);
  nand NAND2_301(g13529,g12611,g3410);
  nand NAND2_302(g13535,g12657,g3566);
  nand NAND2_303(g13536,g12711,g3722);
  nand NAND2_304(g13537,g12565,g3254);
  nand NAND2_305(g13538,g12565,g3254);
  nand NAND2_306(g13539,g12611,g3410);
  nand NAND2_307(g13540,g12657,g3566);
  nand NAND2_308(g13546,g12711,g3722);
  nand NAND2_309(g13547,g12565,g3254);
  nand NAND2_310(g13548,g12611,g3410);
  nand NAND2_311(g13549,g12611,g3410);
  nand NAND2_312(g13550,g12657,g3566);
  nand NAND2_313(g13551,g12711,g3722);
  nand NAND2_314(g13557,g12611,g3410);
  nand NAND2_315(g13558,g12657,g3566);
  nand NAND2_316(g13559,g12657,g3566);
  nand NAND2_317(g13560,g12711,g3722);
  nand NAND2_318(g13561,g12657,g3566);
  nand NAND2_319(g13562,g12711,g3722);
  nand NAND2_320(g13563,g12711,g3722);
  nand NAND2_321(g13564,g12711,g3722);
  nand NAND2_322(g13599,g12886,g3366);
  nand NAND2_323(g13611,g12926,g3522);
  nand NAND2_324(g13621,g12955,g3678);
  nand NAND2_325(g13633,g12984,g3834);
  nand NAND2_326(g13893,g8580,g12463);
  nand NAND3_0(g13915,g8822,g12473,g12463);
  nand NAND2_327(g13934,g8587,g12478);
  nand NAND2_328(g13957,g10730,g12473);
  nand NAND3_1(g13971,g8846,g12490,g12478);
  nand NAND2_329(g13990,g8594,g12495);
  nand NAND2_330(g14027,g10749,g12490);
  nand NAND3_2(g14041,g8873,g12510,g12495);
  nand NAND2_331(g14060,g8605,g12515);
  nand NAND2_332(g14118,g10767,g12510);
  nand NAND3_3(g14132,g8911,g12527,g12515);
  nand NAND2_333(g14233,g10773,g12527);
  nand NAND3_4(g15454,g9232,g9150,g12780);
  nand NAND3_5(g15540,g9310,g9174,g12819);
  nand NAND3_6(g15618,g9391,g9216,g12857);
  nand NAND2_334(g15660,g13401,g12354);
  nand NAND2_335(g15664,g12565,g6314);
  nand NAND3_7(g15694,g9488,g9277,g12898);
  nand NAND2_336(g15718,g13286,g12354);
  nand NAND2_337(g15719,g13401,g12392);
  nand NAND2_338(g15720,g12565,g6232);
  nand NAND2_339(g15721,g12565,g6314);
  nand NAND2_340(g15723,g12611,g6519);
  nand NAND2_341(g15756,g13313,g12354);
  nand NAND2_342(g15757,g11622,g12392);
  nand NAND2_343(g15758,g12565,g6232);
  nand NAND2_344(g15759,g12565,g6314);
  nand NAND2_345(g15760,g12611,g6369);
  nand NAND2_346(g15761,g12611,g6519);
  nand NAND2_347(g15763,g12657,g6783);
  nand NAND2_348(g15782,g13332,g12354);
  nand NAND2_349(g15783,g11643,g12392);
  nand NAND2_350(g15784,g12565,g6232);
  nand NAND2_351(g15785,g12565,g6314);
  nand NAND2_352(g15786,g12611,g6369);
  nand NAND2_353(g15787,g12611,g6519);
  nand NAND2_354(g15788,g12657,g6574);
  nand NAND2_355(g15789,g12657,g6783);
  nand NAND2_356(g15791,g12711,g7085);
  nand NAND2_357(g15803,g13375,g12354);
  nand NAND2_358(g15804,g11660,g12392);
  nand NAND2_359(g15805,g12565,g6232);
  nand NAND2_360(g15806,g12565,g6314);
  nand NAND2_361(g15807,g12611,g6369);
  nand NAND2_362(g15808,g12611,g6519);
  nand NAND2_363(g15809,g12657,g6574);
  nand NAND2_364(g15810,g12657,g6783);
  nand NAND2_365(g15811,g12711,g6838);
  nand NAND2_366(g15812,g12711,g7085);
  nand NAND2_367(II22062,g12999,g12988);
  nand NAND2_368(II22063,g12999,II22062);
  nand NAND2_369(II22064,g12988,II22062);
  nand NAND2_370(g15814,II22063,II22064);
  nand NAND2_371(g15818,g13024,g12354);
  nand NAND2_372(g15819,g13286,g12392);
  nand NAND2_373(g15820,g12565,g6232);
  nand NAND2_374(g15821,g12565,g6314);
  nand NAND2_375(g15822,g12611,g6369);
  nand NAND2_376(g15823,g12611,g6519);
  nand NAND2_377(g15824,g12657,g6574);
  nand NAND2_378(g15825,g12657,g6783);
  nand NAND2_379(g15826,g12711,g6838);
  nand NAND2_380(g15827,g12711,g7085);
  nand NAND2_381(g15830,g13310,g12392);
  nand NAND2_382(g15831,g13313,g12392);
  nand NAND2_383(g15832,g12565,g6232);
  nand NAND2_384(g15833,g12565,g6314);
  nand NAND2_385(g15834,g12611,g6369);
  nand NAND2_386(g15835,g12611,g6519);
  nand NAND2_387(g15836,g12657,g6574);
  nand NAND2_388(g15837,g12657,g6783);
  nand NAND2_389(g15838,g12711,g6838);
  nand NAND2_390(g15839,g12711,g7085);
  nand NAND2_391(g15841,g13331,g12392);
  nand NAND2_392(g15842,g13332,g12392);
  nand NAND2_393(g15843,g12565,g6314);
  nand NAND2_394(g15844,g12565,g6232);
  nand NAND2_395(g15845,g12565,g6314);
  nand NAND2_396(g15846,g12611,g6369);
  nand NAND2_397(g15847,g12611,g6519);
  nand NAND2_398(g15848,g12657,g6574);
  nand NAND2_399(g15849,g12657,g6783);
  nand NAND2_400(g15850,g12711,g6838);
  nand NAND2_401(g15851,g12711,g7085);
  nand NAND2_402(g15853,g13310,g12354);
  nand NAND2_403(g15854,g13353,g12392);
  nand NAND2_404(g15855,g13354,g12392);
  nand NAND2_405(g15856,g12565,g6232);
  nand NAND2_406(g15857,g12565,g6314);
  nand NAND2_407(g15858,g12565,g6232);
  nand NAND2_408(g15866,g12611,g6519);
  nand NAND2_409(g15867,g12611,g6369);
  nand NAND2_410(g15868,g12611,g6519);
  nand NAND2_411(g15869,g12657,g6574);
  nand NAND2_412(g15870,g12657,g6783);
  nand NAND2_413(g15871,g12711,g6838);
  nand NAND2_414(g15872,g12711,g7085);
  nand NAND2_415(g15877,g13374,g12392);
  nand NAND2_416(g15878,g13375,g12392);
  nand NAND2_417(g15879,g12565,g6232);
  nand NAND2_418(g15887,g12611,g6369);
  nand NAND2_419(g15888,g12611,g6519);
  nand NAND2_420(g15889,g12611,g6369);
  nand NAND2_421(g15897,g12657,g6783);
  nand NAND2_422(g15898,g12657,g6574);
  nand NAND2_423(g15899,g12657,g6783);
  nand NAND2_424(g15900,g12711,g6838);
  nand NAND2_425(g15901,g12711,g7085);
  nand NAND2_426(g15903,g13404,g12392);
  nand NAND2_427(g15912,g12611,g6369);
  nand NAND2_428(g15920,g12657,g6574);
  nand NAND2_429(g15921,g12657,g6783);
  nand NAND2_430(g15922,g12657,g6574);
  nand NAND2_431(g15930,g12711,g7085);
  nand NAND2_432(g15931,g12711,g6838);
  nand NAND2_433(g15932,g12711,g7085);
  nand NAND2_434(g15941,g12657,g6574);
  nand NAND2_435(g15949,g12711,g6838);
  nand NAND2_436(g15950,g12711,g7085);
  nand NAND2_437(g15951,g12711,g6838);
  nand NAND2_438(g15970,g12711,g6838);
  nand NAND2_439(g15990,g12886,g6912);
  nand NAND2_440(g15992,g12886,g6678);
  nand NAND2_441(g15993,g12926,g7162);
  nand NAND2_442(g15995,g12926,g6980);
  nand NAND2_443(g15996,g12955,g7358);
  nand NAND2_444(g15999,g12955,g7230);
  nand NAND2_445(g16000,g12984,g7488);
  nand NAND2_446(g16006,g12984,g7426);
  nand NAND2_447(g16085,g12883,g633);
  nand NAND2_448(g16123,g12923,g1319);
  nand NAND2_449(II22282,g2962,g13348);
  nand NAND2_450(II22283,g2962,II22282);
  nand NAND2_451(II22284,g13348,II22282);
  nand NAND2_452(g16132,II22283,II22284);
  nand NAND2_453(g16174,g12952,g2013);
  nand NAND2_454(II22316,g2934,g13370);
  nand NAND2_455(II22317,g2934,II22316);
  nand NAND2_456(II22318,g13370,II22316);
  nand NAND2_457(g16181,II22317,II22318);
  nand NAND2_458(g16233,g12981,g2707);
  nand NAND2_459(g16341,g12377,g12407);
  nand NAND2_460(g16412,g12565,g3254);
  nand NAND2_461(g16439,g13082,g2912);
  nand NAND2_462(g16442,g12565,g3254);
  nand NAND2_463(g16446,g12611,g3410);
  nand NAND2_464(g16463,g13004,g3018);
  nand NAND2_465(g16536,g15873,g2896);
  nand NAND2_466(II22630,g13507,g15978);
  nand NAND2_467(II22631,g13507,II22630);
  nand NAND2_468(II22632,g15978,II22630);
  nand NAND2_469(g16566,II22631,II22632);
  nand NAND2_470(II22705,g13348,g15661);
  nand NAND2_471(II22706,g13348,II22705);
  nand NAND2_472(II22707,g15661,II22705);
  nand NAND2_473(g16662,II22706,II22707);
  nand NAND2_474(II22884,g13370,g15661);
  nand NAND2_475(II22885,g13370,II22884);
  nand NAND2_476(II22886,g15661,II22884);
  nand NAND2_477(g16935,II22885,II22886);
  nand NAND2_478(II22900,g15022,g14000);
  nand NAND2_479(II22901,g15022,II22900);
  nand NAND2_480(II22902,g14000,II22900);
  nand NAND2_481(g16965,II22901,II22902);
  nand NAND2_482(II22917,g15096,g13945);
  nand NAND2_483(II22918,g15096,II22917);
  nand NAND2_484(II22919,g13945,II22917);
  nand NAND2_485(g16985,II22918,II22919);
  nand NAND2_486(II22924,g15118,g14091);
  nand NAND2_487(II22925,g15118,II22924);
  nand NAND2_488(II22926,g14091,II22924);
  nand NAND2_489(g16986,II22925,II22926);
  nand NAND2_490(II22936,g9150,g13906);
  nand NAND2_491(II22937,g9150,II22936);
  nand NAND2_492(II22938,g13906,II22936);
  nand NAND2_493(g16992,II22937,II22938);
  nand NAND2_494(II22945,g15188,g14015);
  nand NAND2_495(II22946,g15188,II22945);
  nand NAND2_496(II22947,g14015,II22945);
  nand NAND2_497(g16995,II22946,II22947);
  nand NAND2_498(II22952,g15210,g14206);
  nand NAND2_499(II22953,g15210,II22952);
  nand NAND2_500(II22954,g14206,II22952);
  nand NAND2_501(g16996,II22953,II22954);
  nand NAND2_502(II22962,g9161,g13885);
  nand NAND2_503(II22963,g9161,II22962);
  nand NAND2_504(II22964,g13885,II22962);
  nand NAND2_505(g17000,II22963,II22964);
  nand NAND2_506(II22972,g9174,g13962);
  nand NAND2_507(II22973,g9174,II22972);
  nand NAND2_508(II22974,g13962,II22972);
  nand NAND2_509(g17016,II22973,II22974);
  nand NAND2_510(II22981,g15274,g14106);
  nand NAND2_511(II22982,g15274,II22981);
  nand NAND2_512(II22983,g14106,II22981);
  nand NAND2_513(g17019,II22982,II22983);
  nand NAND2_514(II22988,g15296,g14321);
  nand NAND2_515(II22989,g15296,II22988);
  nand NAND2_516(II22990,g14321,II22988);
  nand NAND2_517(g17020,II22989,II22990);
  nand NAND2_518(II22998,g9187,g13872);
  nand NAND2_519(II22999,g9187,II22998);
  nand NAND2_520(II23000,g13872,II22998);
  nand NAND2_521(g17024,II22999,II23000);
  nand NAND2_522(II23008,g9203,g13926);
  nand NAND2_523(II23009,g9203,II23008);
  nand NAND2_524(II23010,g13926,II23008);
  nand NAND2_525(g17030,II23009,II23010);
  nand NAND2_526(II23018,g9216,g14032);
  nand NAND2_527(II23019,g9216,II23018);
  nand NAND2_528(II23020,g14032,II23018);
  nand NAND2_529(g17046,II23019,II23020);
  nand NAND2_530(II23027,g15366,g14221);
  nand NAND2_531(II23028,g15366,II23027);
  nand NAND2_532(II23029,g14221,II23027);
  nand NAND2_533(g17049,II23028,II23029);
  nand NAND2_534(II23034,g9232,g13864);
  nand NAND2_535(II23035,g9232,II23034);
  nand NAND2_536(II23036,g13864,II23034);
  nand NAND2_537(g17050,II23035,II23036);
  nand NAND2_538(II23045,g9248,g13894);
  nand NAND2_539(II23046,g9248,II23045);
  nand NAND2_540(II23047,g13894,II23045);
  nand NAND2_541(g17058,II23046,II23047);
  nand NAND2_542(II23055,g9264,g13982);
  nand NAND2_543(II23056,g9264,II23055);
  nand NAND2_544(II23057,g13982,II23055);
  nand NAND2_545(g17064,II23056,II23057);
  nand NAND2_546(II23065,g9277,g14123);
  nand NAND2_547(II23066,g9277,II23065);
  nand NAND2_548(II23067,g14123,II23065);
  nand NAND2_549(g17080,II23066,II23067);
  nand NAND2_550(II23074,g9293,g13856);
  nand NAND2_551(II23075,g9293,II23074);
  nand NAND2_552(II23076,g13856,II23074);
  nand NAND2_553(g17083,II23075,II23076);
  nand NAND2_554(II23082,g9310,g13879);
  nand NAND2_555(II23083,g9310,II23082);
  nand NAND2_556(II23084,g13879,II23082);
  nand NAND2_557(g17085,II23083,II23084);
  nand NAND2_558(II23093,g9326,g13935);
  nand NAND2_559(II23094,g9326,II23093);
  nand NAND2_560(II23095,g13935,II23093);
  nand NAND2_561(g17093,II23094,II23095);
  nand NAND2_562(II23103,g9342,g14052);
  nand NAND2_563(II23104,g9342,II23103);
  nand NAND2_564(II23105,g14052,II23103);
  nand NAND2_565(g17099,II23104,II23105);
  nand NAND2_566(II23113,g9356,g13848);
  nand NAND2_567(II23114,g9356,II23113);
  nand NAND2_568(II23115,g13848,II23113);
  nand NAND2_569(g17115,II23114,II23115);
  nand NAND2_570(g17118,g13915,g13893);
  nand NAND2_571(II23123,g9374,g13866);
  nand NAND2_572(II23124,g9374,II23123);
  nand NAND2_573(II23125,g13866,II23123);
  nand NAND2_574(g17121,II23124,II23125);
  nand NAND2_575(II23131,g9391,g13901);
  nand NAND2_576(II23132,g9391,II23131);
  nand NAND2_577(II23133,g13901,II23131);
  nand NAND2_578(g17123,II23132,II23133);
  nand NAND2_579(II23142,g9407,g13991);
  nand NAND2_580(II23143,g9407,II23142);
  nand NAND2_581(II23144,g13991,II23142);
  nand NAND2_582(g17131,II23143,II23144);
  nand NAND2_583(II23152,g9427,g14061);
  nand NAND2_584(II23153,g9427,II23152);
  nand NAND2_585(II23154,g14061,II23152);
  nand NAND2_586(g17137,II23153,II23154);
  nand NAND2_587(g17139,g13957,g13915);
  nand NAND2_588(II23161,g9453,g13857);
  nand NAND2_589(II23162,g9453,II23161);
  nand NAND2_590(II23163,g13857,II23161);
  nand NAND2_591(g17142,II23162,II23163);
  nand NAND2_592(g17145,g13971,g13934);
  nand NAND2_593(II23171,g9471,g13881);
  nand NAND2_594(II23172,g9471,II23171);
  nand NAND2_595(II23173,g13881,II23171);
  nand NAND2_596(g17148,II23172,II23173);
  nand NAND2_597(II23179,g9488,g13942);
  nand NAND2_598(II23180,g9488,II23179);
  nand NAND2_599(II23181,g13942,II23179);
  nand NAND2_600(g17150,II23180,II23181);
  nand NAND2_601(II23190,g9507,g13999);
  nand NAND2_602(II23191,g9507,II23190);
  nand NAND2_603(II23192,g13999,II23190);
  nand NAND2_604(g17158,II23191,II23192);
  nand NAND2_605(g17159,g14642,g14657);
  nand NAND2_606(II23198,g9569,g14176);
  nand NAND2_607(II23199,g9569,II23198);
  nand NAND2_608(II23200,g14176,II23198);
  nand NAND2_609(g17160,II23199,II23200);
  nand NAND2_610(g17162,g14027,g13971);
  nand NAND2_611(II23207,g9595,g13867);
  nand NAND2_612(II23208,g9595,II23207);
  nand NAND2_613(II23209,g13867,II23207);
  nand NAND2_614(g17165,II23208,II23209);
  nand NAND2_615(g17168,g14041,g13990);
  nand NAND2_616(II23217,g9613,g13903);
  nand NAND2_617(II23218,g9613,II23217);
  nand NAND2_618(II23219,g13903,II23217);
  nand NAND2_619(g17171,II23218,II23219);
  nand NAND2_620(II23225,g9649,g14090);
  nand NAND2_621(II23226,g9649,II23225);
  nand NAND2_622(II23227,g14090,II23225);
  nand NAND2_623(g17173,II23226,II23227);
  nand NAND2_624(g17174,g14669,g14691);
  nand NAND2_625(II23233,g9711,g14291);
  nand NAND2_626(II23234,g9711,II23233);
  nand NAND2_627(II23235,g14291,II23233);
  nand NAND2_628(g17175,II23234,II23235);
  nand NAND2_629(g17177,g14118,g14041);
  nand NAND2_630(II23242,g9737,g13882);
  nand NAND2_631(II23243,g9737,II23242);
  nand NAND2_632(II23244,g13882,II23242);
  nand NAND2_633(g17180,II23243,II23244);
  nand NAND2_634(g17183,g14132,g14060);
  nand NAND2_635(II23256,g9795,g14205);
  nand NAND2_636(II23257,g9795,II23256);
  nand NAND2_637(II23258,g14205,II23256);
  nand NAND2_638(g17190,II23257,II23258);
  nand NAND2_639(g17191,g14703,g14725);
  nand NAND2_640(II23264,g9857,g14413);
  nand NAND2_641(II23265,g9857,II23264);
  nand NAND2_642(II23266,g14413,II23264);
  nand NAND2_643(g17192,II23265,II23266);
  nand NAND2_644(g17194,g14233,g14132);
  nand NAND2_645(II23277,g9941,g14320);
  nand NAND2_646(II23278,g9941,II23277);
  nand NAND2_647(II23279,g14320,II23277);
  nand NAND2_648(g17201,II23278,II23279);
  nand NAND2_649(g17202,g14737,g14753);
  nand NAND2_650(II23806,g14062,g9150);
  nand NAND2_651(II23807,g14062,II23806);
  nand NAND2_652(II23808,g9150,II23806);
  nand NAND2_653(g17729,II23807,II23808);
  nand NAND2_654(II23878,g14001,g9187);
  nand NAND2_655(II23879,g14001,II23878);
  nand NAND2_656(II23880,g9187,II23878);
  nand NAND2_657(g17807,II23879,II23880);
  nand NAND2_658(II23893,g14177,g9174);
  nand NAND2_659(II23894,g14177,II23893);
  nand NAND2_660(II23895,g9174,II23893);
  nand NAND2_661(g17830,II23894,II23895);
  nand NAND2_662(II23941,g13946,g9293);
  nand NAND2_663(II23942,g13946,II23941);
  nand NAND2_664(II23943,g9293,II23941);
  nand NAND2_665(g17887,II23942,II23943);
  nand NAND2_666(II23958,g6513,g14171);
  nand NAND2_667(II23959,g6513,II23958);
  nand NAND2_668(II23960,g14171,II23958);
  nand NAND2_669(g17913,II23959,II23960);
  nand NAND2_670(II23966,g14092,g9248);
  nand NAND2_671(II23967,g14092,II23966);
  nand NAND2_672(II23968,g9248,II23966);
  nand NAND2_673(g17919,II23967,II23968);
  nand NAND2_674(II23981,g14292,g9216);
  nand NAND2_675(II23982,g14292,II23981);
  nand NAND2_676(II23983,g9216,II23981);
  nand NAND2_677(g17942,II23982,II23983);
  nand NAND2_678(II24005,g7548,g15814);
  nand NAND2_679(II24006,g7548,II24005);
  nand NAND2_680(II24007,g15814,II24005);
  nand NAND2_681(g17968,II24006,II24007);
  nand NAND2_682(II24015,g13907,g9427);
  nand NAND2_683(II24016,g13907,II24015);
  nand NAND2_684(II24017,g9427,II24015);
  nand NAND2_685(g17979,II24016,II24017);
  nand NAND2_686(g17985,g14641,g9636);
  nand NAND2_687(II24028,g6201,g14086);
  nand NAND2_688(II24029,g6201,II24028);
  nand NAND2_689(II24030,g14086,II24028);
  nand NAND2_690(g17992,II24029,II24030);
  nand NAND2_691(II24036,g14016,g9374);
  nand NAND2_692(II24037,g14016,II24036);
  nand NAND2_693(II24038,g9374,II24036);
  nand NAND2_694(g17998,II24037,II24038);
  nand NAND2_695(II24053,g6777,g14286);
  nand NAND2_696(II24054,g6777,II24053);
  nand NAND2_697(II24055,g14286,II24053);
  nand NAND2_698(g18024,II24054,II24055);
  nand NAND2_699(II24061,g14207,g9326);
  nand NAND2_700(II24062,g14207,II24061);
  nand NAND2_701(II24063,g9326,II24061);
  nand NAND2_702(g18030,II24062,II24063);
  nand NAND2_703(II24076,g14414,g9277);
  nand NAND2_704(II24077,g14414,II24076);
  nand NAND2_705(II24078,g9277,II24076);
  nand NAND2_706(g18053,II24077,II24078);
  nand NAND2_707(II24091,g13886,g15096);
  nand NAND2_708(II24092,g13886,II24091);
  nand NAND2_709(II24093,g15096,II24091);
  nand NAND2_710(g18079,II24092,II24093);
  nand NAND2_711(II24102,g6363,g14011);
  nand NAND2_712(II24103,g6363,II24102);
  nand NAND2_713(II24104,g14011,II24102);
  nand NAND2_714(g18090,II24103,II24104);
  nand NAND2_715(II24110,g13963,g9569);
  nand NAND2_716(II24111,g13963,II24110);
  nand NAND2_717(II24112,g9569,II24110);
  nand NAND2_718(g18096,II24111,II24112);
  nand NAND2_719(g18102,g14668,g9782);
  nand NAND2_720(II24123,g6290,g14201);
  nand NAND2_721(II24124,g6290,II24123);
  nand NAND2_722(II24125,g14201,II24123);
  nand NAND2_723(g18109,II24124,II24125);
  nand NAND2_724(II24131,g14107,g9471);
  nand NAND2_725(II24132,g14107,II24131);
  nand NAND2_726(II24133,g9471,II24131);
  nand NAND2_727(g18115,II24132,II24133);
  nand NAND2_728(II24148,g7079,g14408);
  nand NAND2_729(II24149,g7079,II24148);
  nand NAND2_730(II24150,g14408,II24148);
  nand NAND2_731(g18141,II24149,II24150);
  nand NAND2_732(II24156,g14322,g9407);
  nand NAND2_733(II24157,g14322,II24156);
  nand NAND2_734(II24158,g9407,II24156);
  nand NAND2_735(g18147,II24157,II24158);
  nand NAND2_736(II24178,g13873,g9161);
  nand NAND2_737(II24179,g13873,II24178);
  nand NAND2_738(II24180,g9161,II24178);
  nand NAND2_739(g18183,II24179,II24180);
  nand NAND2_740(II24186,g6177,g13958);
  nand NAND2_741(II24187,g6177,II24186);
  nand NAND2_742(II24188,g13958,II24186);
  nand NAND2_743(g18189,II24187,II24188);
  nand NAND2_744(II24194,g13927,g15188);
  nand NAND2_745(II24195,g13927,II24194);
  nand NAND2_746(II24196,g15188,II24194);
  nand NAND2_747(g18195,II24195,II24196);
  nand NAND2_748(II24205,g6568,g14102);
  nand NAND2_749(II24206,g6568,II24205);
  nand NAND2_750(II24207,g14102,II24205);
  nand NAND2_751(g18206,II24206,II24207);
  nand NAND2_752(II24213,g14033,g9711);
  nand NAND2_753(II24214,g14033,II24213);
  nand NAND2_754(II24215,g9711,II24213);
  nand NAND2_755(g18212,II24214,II24215);
  nand NAND2_756(g18218,g14702,g9928);
  nand NAND2_757(II24226,g6427,g14316);
  nand NAND2_758(II24227,g6427,II24226);
  nand NAND2_759(II24228,g14316,II24226);
  nand NAND2_760(g18225,II24227,II24228);
  nand NAND2_761(II24234,g14222,g9613);
  nand NAND2_762(II24235,g14222,II24234);
  nand NAND2_763(II24236,g9613,II24234);
  nand NAND2_764(g18231,II24235,II24236);
  nand NAND2_765(II24251,g7329,g14520);
  nand NAND2_766(II24252,g7329,II24251);
  nand NAND2_767(II24253,g14520,II24251);
  nand NAND2_768(g18257,II24252,II24253);
  nand NAND2_769(II24263,g14342,g9232);
  nand NAND2_770(II24264,g14342,II24263);
  nand NAND2_771(II24265,g9232,II24263);
  nand NAND2_772(g18270,II24264,II24265);
  nand NAND2_773(II24271,g6180,g13922);
  nand NAND2_774(II24272,g6180,II24271);
  nand NAND2_775(II24273,g13922,II24271);
  nand NAND2_776(g18276,II24272,II24273);
  nand NAND2_777(II24278,g6284,g13918);
  nand NAND2_778(II24279,g6284,II24278);
  nand NAND2_779(II24280,g13918,II24278);
  nand NAND2_780(g18277,II24279,II24280);
  nand NAND2_781(II24290,g13895,g9203);
  nand NAND2_782(II24291,g13895,II24290);
  nand NAND2_783(II24292,g9203,II24290);
  nand NAND2_784(g18290,II24291,II24292);
  nand NAND2_785(II24298,g6209,g14028);
  nand NAND2_786(II24299,g6209,II24298);
  nand NAND2_787(II24300,g14028,II24298);
  nand NAND2_788(g18296,II24299,II24300);
  nand NAND2_789(II24306,g13983,g15274);
  nand NAND2_790(II24307,g13983,II24306);
  nand NAND2_791(II24308,g15274,II24306);
  nand NAND2_792(g18302,II24307,II24308);
  nand NAND2_793(II24317,g6832,g14217);
  nand NAND2_794(II24318,g6832,II24317);
  nand NAND2_795(II24319,g14217,II24317);
  nand NAND2_796(g18313,II24318,II24319);
  nand NAND2_797(II24325,g14124,g9857);
  nand NAND2_798(II24326,g14124,II24325);
  nand NAND2_799(II24327,g9857,II24325);
  nand NAND2_800(g18319,II24326,II24327);
  nand NAND2_801(g18325,g14736,g10082);
  nand NAND2_802(II24338,g6632,g14438);
  nand NAND2_803(II24339,g6632,II24338);
  nand NAND2_804(II24340,g14438,II24338);
  nand NAND2_805(g18332,II24339,II24340);
  nand NAND2_806(II24351,g14238,g9356);
  nand NAND2_807(II24352,g14238,II24351);
  nand NAND2_808(II24353,g9356,II24351);
  nand NAND2_809(g18346,II24352,II24353);
  nand NAND2_810(II24361,g6157,g14525);
  nand NAND2_811(II24362,g6157,II24361);
  nand NAND2_812(II24363,g14525,II24361);
  nand NAND2_813(g18354,II24362,II24363);
  nand NAND2_814(II24372,g14454,g9310);
  nand NAND2_815(II24373,g14454,II24372);
  nand NAND2_816(II24374,g9310,II24372);
  nand NAND2_817(g18363,II24373,II24374);
  nand NAND2_818(II24380,g6212,g13978);
  nand NAND2_819(II24381,g6212,II24380);
  nand NAND2_820(II24382,g13978,II24380);
  nand NAND2_821(g18369,II24381,II24382);
  nand NAND2_822(II24387,g6421,g13974);
  nand NAND2_823(II24388,g6421,II24387);
  nand NAND2_824(II24389,g13974,II24387);
  nand NAND2_825(g18370,II24388,II24389);
  nand NAND2_826(II24399,g13936,g9264);
  nand NAND2_827(II24400,g13936,II24399);
  nand NAND2_828(II24401,g9264,II24399);
  nand NAND2_829(g18383,II24400,II24401);
  nand NAND2_830(II24407,g6298,g14119);
  nand NAND2_831(II24408,g6298,II24407);
  nand NAND2_832(II24409,g14119,II24407);
  nand NAND2_833(g18389,II24408,II24409);
  nand NAND2_834(II24415,g14053,g15366);
  nand NAND2_835(II24416,g14053,II24415);
  nand NAND2_836(II24417,g15366,II24415);
  nand NAND2_837(g18395,II24416,II24417);
  nand NAND2_838(II24426,g7134,g14332);
  nand NAND2_839(II24427,g7134,II24426);
  nand NAND2_840(II24428,g14332,II24426);
  nand NAND2_841(g18406,II24427,II24428);
  nand NAND2_842(II24436,g14153,g15022);
  nand NAND2_843(II24437,g14153,II24436);
  nand NAND2_844(II24438,g15022,II24436);
  nand NAND2_845(g18419,II24437,II24438);
  nand NAND2_846(II24443,g14148,g9507);
  nand NAND2_847(II24444,g14148,II24443);
  nand NAND2_848(II24445,g9507,II24443);
  nand NAND2_849(g18424,II24444,II24445);
  nand NAND2_850(II24452,g6142,g14450);
  nand NAND2_851(II24453,g6142,II24452);
  nand NAND2_852(II24454,g14450,II24452);
  nand NAND2_853(g18431,II24453,II24454);
  nand NAND2_854(II24464,g14360,g9453);
  nand NAND2_855(II24465,g14360,II24464);
  nand NAND2_856(II24466,g9453,II24464);
  nand NAND2_857(g18441,II24465,II24466);
  nand NAND2_858(II24474,g6184,g14580);
  nand NAND2_859(II24475,g6184,II24474);
  nand NAND2_860(II24476,g14580,II24474);
  nand NAND2_861(g18449,II24475,II24476);
  nand NAND2_862(II24485,g14541,g9391);
  nand NAND2_863(II24486,g14541,II24485);
  nand NAND2_864(II24487,g9391,II24485);
  nand NAND2_865(g18458,II24486,II24487);
  nand NAND2_866(II24493,g6301,g14048);
  nand NAND2_867(II24494,g6301,II24493);
  nand NAND2_868(II24495,g14048,II24493);
  nand NAND2_869(g18464,II24494,II24495);
  nand NAND2_870(II24500,g6626,g14044);
  nand NAND2_871(II24501,g6626,II24500);
  nand NAND2_872(II24502,g14044,II24500);
  nand NAND2_873(g18465,II24501,II24502);
  nand NAND2_874(II24512,g13992,g9342);
  nand NAND2_875(II24513,g13992,II24512);
  nand NAND2_876(II24514,g9342,II24512);
  nand NAND2_877(g18478,II24513,II24514);
  nand NAND2_878(II24520,g6435,g14234);
  nand NAND2_879(II24521,g6435,II24520);
  nand NAND2_880(II24522,g14234,II24520);
  nand NAND2_881(g18484,II24521,II24522);
  nand NAND2_882(II24530,g6707,g14355);
  nand NAND2_883(II24531,g6707,II24530);
  nand NAND2_884(II24532,g14355,II24530);
  nand NAND2_885(g18491,II24531,II24532);
  nand NAND2_886(II24537,g14268,g15118);
  nand NAND2_887(II24538,g14268,II24537);
  nand NAND2_888(II24539,g15118,II24537);
  nand NAND2_889(g18492,II24538,II24539);
  nand NAND2_890(II24544,g14263,g9649);
  nand NAND2_891(II24545,g14263,II24544);
  nand NAND2_892(II24546,g9649,II24544);
  nand NAND2_893(g18497,II24545,II24546);
  nand NAND2_894(II24553,g6163,g14537);
  nand NAND2_895(II24554,g6163,II24553);
  nand NAND2_896(II24555,g14537,II24553);
  nand NAND2_897(g18504,II24554,II24555);
  nand NAND2_898(II24565,g14472,g9595);
  nand NAND2_899(II24566,g14472,II24565);
  nand NAND2_900(II24567,g9595,II24565);
  nand NAND2_901(g18514,II24566,II24567);
  nand NAND2_902(II24575,g6216,g14614);
  nand NAND2_903(II24576,g6216,II24575);
  nand NAND2_904(II24577,g14614,II24575);
  nand NAND2_905(g18522,II24576,II24577);
  nand NAND2_906(II24586,g14596,g9488);
  nand NAND2_907(II24587,g14596,II24586);
  nand NAND2_908(II24588,g9488,II24586);
  nand NAND2_909(g18531,II24587,II24588);
  nand NAND2_910(II24594,g6438,g14139);
  nand NAND2_911(II24595,g6438,II24594);
  nand NAND2_912(II24596,g14139,II24594);
  nand NAND2_913(g18537,II24595,II24596);
  nand NAND2_914(II24601,g6890,g14135);
  nand NAND2_915(II24602,g6890,II24601);
  nand NAND2_916(II24603,g14135,II24601);
  nand NAND2_917(g18538,II24602,II24603);
  nand NAND2_918(II24611,g15814,g15978);
  nand NAND2_919(II24612,g15814,II24611);
  nand NAND2_920(II24613,g15978,II24611);
  nand NAND2_921(g18542,II24612,II24613);
  nand NAND2_922(II24624,g6136,g14252);
  nand NAND2_923(II24625,g6136,II24624);
  nand NAND2_924(II24626,g14252,II24624);
  nand NAND2_925(g18553,II24625,II24626);
  nand NAND2_926(II24632,g7009,g14467);
  nand NAND2_927(II24633,g7009,II24632);
  nand NAND2_928(II24634,g14467,II24632);
  nand NAND2_929(g18555,II24633,II24634);
  nand NAND2_930(II24639,g14390,g15210);
  nand NAND2_931(II24640,g14390,II24639);
  nand NAND2_932(II24641,g15210,II24639);
  nand NAND2_933(g18556,II24640,II24641);
  nand NAND2_934(II24646,g14385,g9795);
  nand NAND2_935(II24647,g14385,II24646);
  nand NAND2_936(II24648,g9795,II24646);
  nand NAND2_937(g18561,II24647,II24648);
  nand NAND2_938(II24655,g6190,g14592);
  nand NAND2_939(II24656,g6190,II24655);
  nand NAND2_940(II24657,g14592,II24655);
  nand NAND2_941(g18568,II24656,II24657);
  nand NAND2_942(II24667,g14559,g9737);
  nand NAND2_943(II24668,g14559,II24667);
  nand NAND2_944(II24669,g9737,II24667);
  nand NAND2_945(g18578,II24668,II24669);
  nand NAND2_946(II24677,g6305,g14637);
  nand NAND2_947(II24678,g6305,II24677);
  nand NAND2_948(II24679,g14637,II24677);
  nand NAND2_949(g18586,II24678,II24679);
  nand NAND2_950(II24694,g6146,g14374);
  nand NAND2_951(II24695,g6146,II24694);
  nand NAND2_952(II24696,g14374,II24694);
  nand NAND2_953(g18603,II24695,II24696);
  nand NAND2_954(II24702,g7259,g14554);
  nand NAND2_955(II24703,g7259,II24702);
  nand NAND2_956(II24704,g14554,II24702);
  nand NAND2_957(g18605,II24703,II24704);
  nand NAND2_958(II24709,g14502,g15296);
  nand NAND2_959(II24710,g14502,II24709);
  nand NAND2_960(II24711,g15296,II24709);
  nand NAND2_961(g18606,II24710,II24711);
  nand NAND2_962(II24716,g14497,g9941);
  nand NAND2_963(II24717,g14497,II24716);
  nand NAND2_964(II24718,g9941,II24716);
  nand NAND2_965(g18611,II24717,II24718);
  nand NAND2_966(II24725,g6222,g14626);
  nand NAND2_967(II24726,g6222,II24725);
  nand NAND2_968(II24727,g14626,II24725);
  nand NAND2_969(g18618,II24726,II24727);
  nand NAND2_970(II24743,g6167,g14486);
  nand NAND2_971(II24744,g6167,II24743);
  nand NAND2_972(II24745,g14486,II24743);
  nand NAND2_973(g18635,II24744,II24745);
  nand NAND2_974(II24751,g7455,g14609);
  nand NAND2_975(II24752,g7455,II24751);
  nand NAND2_976(II24753,g14609,II24751);
  nand NAND2_977(g18637,II24752,II24753);
  nand NAND2_978(II24763,g6194,g14573);
  nand NAND2_979(II24764,g6194,II24763);
  nand NAND2_980(II24765,g14573,II24763);
  nand NAND2_981(g18644,II24764,II24765);
  nand NAND2_982(g18977,g15797,g3006);
  nand NAND2_983(II25030,g8029,g13507);
  nand NAND2_984(II25031,g8029,II25030);
  nand NAND2_985(II25032,g13507,II25030);
  nand NAND2_986(g18980,II25031,II25032);
  nand NAND2_987(g19067,g16554,g16578);
  nand NAND2_988(g19084,g16586,g16602);
  nand NAND2_989(g19103,g18590,g2924);
  nand NAND2_990(g19121,g16682,g16697);
  nand NAND2_991(g19128,g16708,g16728);
  nand NAND2_992(g19135,g16739,g16770);
  nand NAND2_993(g19138,g16781,g16797);
  nand NAND2_994(g19141,g3088,g16825);
  nand NAND2_995(g19152,g5378,g18884);
  nand NAND2_996(II25532,g52,g18179);
  nand NAND2_997(II25533,g52,II25532);
  nand NAND2_998(II25534,g18179,II25532);
  nand NAND2_999(g19261,II25533,II25534);
  nand NAND2_1000(II25539,g92,g18174);
  nand NAND2_1001(II25540,g92,II25539);
  nand NAND2_1002(II25541,g18174,II25539);
  nand NAND2_1003(g19262,II25540,II25541);
  nand NAND2_1004(II25560,g56,g17724);
  nand NAND2_1005(II25561,g56,II25560);
  nand NAND2_1006(II25562,g17724,II25560);
  nand NAND2_1007(g19271,II25561,II25562);
  nand NAND2_1008(II25571,g740,g18286);
  nand NAND2_1009(II25572,g740,II25571);
  nand NAND2_1010(II25573,g18286,II25571);
  nand NAND2_1011(g19276,II25572,II25573);
  nand NAND2_1012(II25578,g780,g18281);
  nand NAND2_1013(II25579,g780,II25578);
  nand NAND2_1014(II25580,g18281,II25578);
  nand NAND2_1015(g19277,II25579,II25580);
  nand NAND2_1016(II25595,g61,g18074);
  nand NAND2_1017(II25596,g61,II25595);
  nand NAND2_1018(II25597,g18074,II25595);
  nand NAND2_1019(g19286,II25596,II25597);
  nand NAND3_8(g19288,g14685,g8580,g17057);
  nand NAND2_1020(II25605,g744,g17825);
  nand NAND2_1021(II25606,g744,II25605);
  nand NAND2_1022(II25607,g17825,II25605);
  nand NAND2_1023(g19290,II25606,II25607);
  nand NAND2_1024(II25616,g1426,g18379);
  nand NAND2_1025(II25617,g1426,II25616);
  nand NAND2_1026(II25618,g18379,II25616);
  nand NAND2_1027(g19295,II25617,II25618);
  nand NAND2_1028(II25623,g1466,g18374);
  nand NAND2_1029(II25624,g1466,II25623);
  nand NAND2_1030(II25625,g18374,II25623);
  nand NAND2_1031(g19296,II25624,II25625);
  nand NAND2_1032(II25633,g65,g17640);
  nand NAND2_1033(II25634,g65,II25633);
  nand NAND2_1034(II25635,g17640,II25633);
  nand NAND2_1035(g19300,II25634,II25635);
  nand NAND2_1036(II25643,g749,g18190);
  nand NAND2_1037(II25644,g749,II25643);
  nand NAND2_1038(II25645,g18190,II25643);
  nand NAND2_1039(g19304,II25644,II25645);
  nand NAND3_9(g19306,g14719,g8587,g17092);
  nand NAND2_1040(II25653,g1430,g17937);
  nand NAND2_1041(II25654,g1430,II25653);
  nand NAND2_1042(II25655,g17937,II25653);
  nand NAND2_1043(g19308,II25654,II25655);
  nand NAND2_1044(II25664,g2120,g18474);
  nand NAND2_1045(II25665,g2120,II25664);
  nand NAND2_1046(II25666,g18474,II25664);
  nand NAND2_1047(g19313,II25665,II25666);
  nand NAND2_1048(II25671,g2160,g18469);
  nand NAND2_1049(II25672,g2160,II25671);
  nand NAND2_1050(II25673,g18469,II25671);
  nand NAND2_1051(g19314,II25672,II25673);
  nand NAND2_1052(II25681,g70,g17974);
  nand NAND2_1053(II25682,g70,II25681);
  nand NAND2_1054(II25683,g17974,II25681);
  nand NAND2_1055(g19318,II25682,II25683);
  nand NAND2_1056(II25690,g753,g17741);
  nand NAND2_1057(II25691,g753,II25690);
  nand NAND2_1058(II25692,g17741,II25690);
  nand NAND2_1059(g19321,II25691,II25692);
  nand NAND2_1060(II25700,g1435,g18297);
  nand NAND2_1061(II25701,g1435,II25700);
  nand NAND2_1062(II25702,g18297,II25700);
  nand NAND2_1063(g19325,II25701,II25702);
  nand NAND3_10(g19327,g14747,g8594,g17130);
  nand NAND2_1064(II25710,g2124,g18048);
  nand NAND2_1065(II25711,g2124,II25710);
  nand NAND2_1066(II25712,g18048,II25710);
  nand NAND2_1067(g19329,II25711,II25712);
  nand NAND2_1068(II25721,g74,g18341);
  nand NAND2_1069(II25722,g74,II25721);
  nand NAND2_1070(II25723,g18341,II25721);
  nand NAND2_1071(g19334,II25722,II25723);
  nand NAND2_1072(II25731,g758,g18091);
  nand NAND2_1073(II25732,g758,II25731);
  nand NAND2_1074(II25733,g18091,II25731);
  nand NAND2_1075(g19345,II25732,II25733);
  nand NAND2_1076(II25740,g1439,g17842);
  nand NAND2_1077(II25741,g1439,II25740);
  nand NAND2_1078(II25742,g17842,II25740);
  nand NAND2_1079(g19348,II25741,II25742);
  nand NAND2_1080(II25750,g2129,g18390);
  nand NAND2_1081(II25751,g2129,II25750);
  nand NAND2_1082(II25752,g18390,II25750);
  nand NAND2_1083(g19352,II25751,II25752);
  nand NAND3_11(g19354,g14768,g8605,g17157);
  nand NAND2_1084(II25761,g79,g17882);
  nand NAND2_1085(II25762,g79,II25761);
  nand NAND2_1086(II25763,g17882,II25761);
  nand NAND2_1087(g19357,II25762,II25763);
  nand NAND2_1088(II25771,g762,g18436);
  nand NAND2_1089(II25772,g762,II25771);
  nand NAND2_1090(II25773,g18436,II25771);
  nand NAND2_1091(g19368,II25772,II25773);
  nand NAND2_1092(II25781,g1444,g18207);
  nand NAND2_1093(II25782,g1444,II25781);
  nand NAND2_1094(II25783,g18207,II25781);
  nand NAND2_1095(g19379,II25782,II25783);
  nand NAND2_1096(II25790,g2133,g17954);
  nand NAND2_1097(II25791,g2133,II25790);
  nand NAND2_1098(II25792,g17954,II25790);
  nand NAND2_1099(g19382,II25791,II25792);
  nand NAND2_1100(II25800,g83,g18265);
  nand NAND2_1101(II25801,g83,II25800);
  nand NAND2_1102(II25802,g18265,II25800);
  nand NAND2_1103(g19386,II25801,II25802);
  nand NAND2_1104(II25809,g767,g17993);
  nand NAND2_1105(II25810,g767,II25809);
  nand NAND2_1106(II25811,g17993,II25809);
  nand NAND2_1107(g19389,II25810,II25811);
  nand NAND2_1108(II25819,g1448,g18509);
  nand NAND2_1109(II25820,g1448,II25819);
  nand NAND2_1110(II25821,g18509,II25819);
  nand NAND2_1111(g19400,II25820,II25821);
  nand NAND2_1112(II25829,g2138,g18314);
  nand NAND2_1113(II25830,g2138,II25829);
  nand NAND2_1114(II25831,g18314,II25829);
  nand NAND2_1115(g19411,II25830,II25831);
  nand NAND2_1116(II25838,g88,g17802);
  nand NAND2_1117(II25839,g88,II25838);
  nand NAND2_1118(II25840,g17802,II25838);
  nand NAND2_1119(g19414,II25839,II25840);
  nand NAND2_1120(II25846,g771,g18358);
  nand NAND2_1121(II25847,g771,II25846);
  nand NAND2_1122(II25848,g18358,II25846);
  nand NAND2_1123(g19416,II25847,II25848);
  nand NAND2_1124(II25855,g1453,g18110);
  nand NAND2_1125(II25856,g1453,II25855);
  nand NAND2_1126(II25857,g18110,II25855);
  nand NAND2_1127(g19419,II25856,II25857);
  nand NAND2_1128(II25865,g2142,g18573);
  nand NAND2_1129(II25866,g2142,II25865);
  nand NAND2_1130(II25867,g18573,II25865);
  nand NAND2_1131(g19430,II25866,II25867);
  nand NAND2_1132(II25880,g776,g17914);
  nand NAND2_1133(II25881,g776,II25880);
  nand NAND2_1134(II25882,g17914,II25880);
  nand NAND2_1135(g19451,II25881,II25882);
  nand NAND2_1136(II25888,g1457,g18453);
  nand NAND2_1137(II25889,g1457,II25888);
  nand NAND2_1138(II25890,g18453,II25888);
  nand NAND2_1139(g19453,II25889,II25890);
  nand NAND2_1140(II25897,g2147,g18226);
  nand NAND2_1141(II25898,g2147,II25897);
  nand NAND2_1142(II25899,g18226,II25897);
  nand NAND2_1143(g19456,II25898,II25899);
  nand NAND2_1144(II25913,g1462,g18025);
  nand NAND2_1145(II25914,g1462,II25913);
  nand NAND2_1146(II25915,g18025,II25913);
  nand NAND2_1147(g19478,II25914,II25915);
  nand NAND2_1148(II25921,g2151,g18526);
  nand NAND2_1149(II25922,g2151,II25921);
  nand NAND2_1150(II25923,g18526,II25921);
  nand NAND2_1151(g19480,II25922,II25923);
  nand NAND2_1152(II25938,g2156,g18142);
  nand NAND2_1153(II25939,g2156,II25938);
  nand NAND2_1154(II25940,g18142,II25938);
  nand NAND2_1155(g19501,II25939,II25940);
  nand NAND2_1156(g19865,g16607,g9636);
  nand NAND2_1157(g19896,g16625,g9782);
  nand NAND2_1158(g19921,g16639,g9928);
  nand NAND2_1159(g19936,g16650,g10082);
  nand NAND2_1160(g19954,g17186,g92);
  nand NAND2_1161(g19984,g17197,g780);
  nand NAND2_1162(g20022,g17204,g1466);
  nand NAND2_1163(g20064,g17209,g2160);
  nand NAND2_1164(g20473,g18085,g646);
  nand NAND2_1165(g20481,g18201,g1332);
  nand NAND2_1166(g20487,g18308,g2026);
  nand NAND2_1167(g20493,g18401,g2720);
  nand NAND2_1168(g20497,g5410,g18886);
  nand NAND2_1169(g20522,g16501,g16515);
  nand NAND2_1170(g20537,g18626,g3036);
  nand NAND2_1171(g20542,g16523,g16546);
  nand NAND2_1172(g20633,g20164,g3254);
  nand NAND2_1173(g20648,g20164,g3254);
  nand NAND2_1174(g20658,g20198,g3410);
  nand NAND2_1175(g20672,g20164,g3254);
  nand NAND2_1176(g20683,g20198,g3410);
  nand NAND2_1177(g20693,g20228,g3566);
  nand NAND2_1178(g20700,g20153,g2903);
  nand NAND2_1179(g20703,g20164,g3254);
  nand NAND2_1180(g20707,g20198,g3410);
  nand NAND2_1181(g20718,g20228,g3566);
  nand NAND2_1182(g20728,g20255,g3722);
  nand NAND2_1183(g20738,g20198,g3410);
  nand NAND2_1184(g20742,g20228,g3566);
  nand NAND2_1185(g20753,g20255,g3722);
  nand NAND2_1186(g20775,g20228,g3566);
  nand NAND2_1187(g20779,g20255,g3722);
  nand NAND2_1188(g20805,g20255,g3722);
  nand NAND2_1189(g20825,g19219,g15959);
  nand NAND2_1190(g21659,g20164,g6314);
  nand NAND2_1191(II28189,g14079,g19444);
  nand NAND2_1192(II28190,g14079,II28189);
  nand NAND2_1193(II28191,g19444,II28189);
  nand NAND2_1194(g21660,II28190,II28191);
  nand NAND2_1195(g21685,g20164,g6232);
  nand NAND2_1196(g21686,g20164,g6314);
  nand NAND2_1197(g21688,g20198,g6519);
  nand NAND2_1198(II28217,g14194,g19471);
  nand NAND2_1199(II28218,g14194,II28217);
  nand NAND2_1200(II28219,g19471,II28217);
  nand NAND2_1201(g21689,II28218,II28219);
  nand NAND2_1202(g21714,g20164,g6232);
  nand NAND2_1203(g21715,g20164,g6314);
  nand NAND4_1(g21720,g14256,g15177,g19871,g19842);
  nand NAND2_1204(g21721,g20198,g6369);
  nand NAND2_1205(g21722,g20198,g6519);
  nand NAND2_1206(g21724,g20228,g6783);
  nand NAND2_1207(II28247,g14309,g19494);
  nand NAND2_1208(II28248,g14309,II28247);
  nand NAND2_1209(II28249,g19494,II28247);
  nand NAND2_1210(g21725,II28248,II28249);
  nand NAND2_1211(g21736,g20164,g6232);
  nand NAND2_1212(g21737,g20164,g6314);
  nand NAND2_1213(g21740,g20198,g6369);
  nand NAND2_1214(g21741,g20198,g6519);
  nand NAND4_2(g21746,g14378,g15263,g19902,g19875);
  nand NAND2_1215(g21747,g20228,g6574);
  nand NAND2_1216(g21748,g20228,g6783);
  nand NAND2_1217(g21750,g20255,g7085);
  nand NAND2_1218(II28271,g14431,g19515);
  nand NAND2_1219(II28272,g14431,II28271);
  nand NAND2_1220(II28273,g19515,II28271);
  nand NAND2_1221(g21751,II28272,II28273);
  nand NAND2_1222(g21759,g20164,g6232);
  nand NAND2_1223(g21760,g20198,g6369);
  nand NAND2_1224(g21761,g20198,g6519);
  nand NAND2_1225(g21764,g20228,g6574);
  nand NAND2_1226(g21765,g20228,g6783);
  nand NAND4_3(g21770,g14490,g15355,g19927,g19906);
  nand NAND2_1227(g21771,g20255,g6838);
  nand NAND2_1228(g21772,g20255,g7085);
  nand NAND2_1229(g21775,g20198,g6369);
  nand NAND2_1230(g21776,g20228,g6574);
  nand NAND2_1231(g21777,g20228,g6783);
  nand NAND2_1232(g21780,g20255,g6838);
  nand NAND2_1233(g21781,g20255,g7085);
  nand NAND4_4(g21786,g14577,g15441,g19942,g19931);
  nand NAND2_1234(g21790,g20228,g6574);
  nand NAND2_1235(g21791,g20255,g6838);
  nand NAND2_1236(g21792,g20255,g7085);
  nand NAND2_1237(g21804,g20255,g6838);
  nand NAND3_12(g21848,g17807,g19181,g19186);
  nand NAND3_13(g21850,g17979,g19187,g19191);
  nand NAND3_14(g21855,g17919,g19188,g19193);
  nand NAND3_15(g21857,g18079,g19192,g19200);
  nand NAND3_16(g21858,g18096,g19194,g19202);
  nand NAND3_17(g21859,g18030,g19195,g19204);
  nand NAND3_18(g21860,g18270,g19201,g19209);
  nand NAND3_19(g21862,g18195,g19203,g19211);
  nand NAND3_20(g21863,g18212,g19205,g19213);
  nand NAND3_21(g21864,g18147,g19206,g19215);
  nand NAND3_22(g21865,g18424,g19210,g19221);
  nand NAND3_23(g21866,g18363,g19212,g19222);
  nand NAND3_24(g21868,g18302,g19214,g19224);
  nand NAND3_25(g21869,g18319,g19216,g19226);
  nand NAND3_26(g21870,g18497,g19223,g19231);
  nand NAND3_27(g21871,g18458,g19225,g19232);
  nand NAND3_28(g21873,g18395,g19227,g19234);
  nand NAND3_29(g21874,g18561,g19233,g19244);
  nand NAND3_30(g21875,g18531,g19235,g19245);
  nand NAND3_31(g21877,g18611,g19246,g19257);
  nand NAND3_32(g21879,g18419,g19250,g19263);
  nand NAND3_33(g21881,g18492,g19264,g19278);
  nand NAND3_34(g21885,g18556,g19279,g19297);
  nand NAND3_35(g21888,g18606,g19298,g19315);
  nand NAND2_1238(g21903,g20008,g3013);
  nand NAND3_36(g21976,g19242,g21120,g19275);
  nand NAND3_37(g21983,g19255,g21139,g19294);
  nand NAND2_1239(g21989,g21048,g18623);
  nand NAND2_1240(g21991,g21501,g21536);
  nand NAND3_38(g21996,g19268,g21159,g19312);
  nand NAND2_1241(g22002,g21065,g21711);
  nand NAND2_1242(g22005,g21540,g21572);
  nand NAND3_39(g22009,g19283,g21179,g19333);
  nand NAND2_1243(g22016,g21576,g21605);
  nand NAND2_1244(g22021,g21609,g21634);
  nand NAND3_40(g22050,g19450,g21244,g19503);
  nand NAND3_41(g22069,g19477,g21253,g19522);
  nand NAND2_1245(g22083,g21774,g21787);
  nand NAND3_42(g22093,g19500,g21261,g19532);
  nand NAND2_1246(g22108,g21789,g21801);
  nand NAND3_43(g22118,g19521,g21269,g19542);
  nand NAND2_1247(g22134,g21803,g21809);
  nand NAND2_1248(g22157,g21811,g21816);
  nand NAND2_1249(II28726,g21887,g13519);
  nand NAND2_1250(II28727,g21887,II28726);
  nand NAND2_1251(II28728,g13519,II28726);
  nand NAND2_1252(g22188,II28727,II28728);
  nand NAND2_1253(II28741,g21890,g13530);
  nand NAND2_1254(II28742,g21890,II28741);
  nand NAND2_1255(II28743,g13530,II28741);
  nand NAND2_1256(g22197,II28742,II28743);
  nand NAND2_1257(II28753,g21893,g13541);
  nand NAND2_1258(II28754,g21893,II28753);
  nand NAND2_1259(II28755,g13541,II28753);
  nand NAND2_1260(g22203,II28754,II28755);
  nand NAND2_1261(II28765,g21901,g13552);
  nand NAND2_1262(II28766,g21901,II28765);
  nand NAND2_1263(II28767,g13552,II28765);
  nand NAND2_1264(g22209,II28766,II28767);
  nand NAND3_44(g22317,g21152,g21241,g21136);
  nand NAND3_45(g22339,g14442,g21149,g10694);
  nand NAND3_46(g22342,g21172,g21249,g21156);
  nand NAND3_47(g22362,g14529,g21169,g10714);
  nand NAND3_48(g22365,g21192,g21258,g21176);
  nand NAND3_49(g22381,g21211,g14442,g10694);
  nand NAND3_50(g22382,g14584,g21189,g10735);
  nand NAND3_51(g22385,g21207,g21266,g21196);
  nand NAND3_52(g22396,g21219,g14529,g10714);
  nand NAND3_53(g22397,g14618,g21204,g10754);
  nand NAND3_54(g22399,g21230,g14584,g10735);
  nand NAND3_55(g22400,g21235,g14618,g10754);
  nand NAND2_1265(g22608,g20842,g20885);
  nand NAND2_1266(g22644,g20850,g20904);
  nand NAND2_1267(g22668,g16075,g21271);
  nand NAND2_1268(g22680,g20858,g20928);
  nand NAND2_1269(g22708,g16113,g21278);
  nand NAND2_1270(g22720,g20866,g20956);
  nand NAND2_1271(g22739,g16164,g21285);
  nand NAND2_1272(g22771,g16223,g21293);
  nand NAND3_56(g22809,g21850,g21848,g21879);
  nand NAND3_57(g22844,g21865,g21860,g21857);
  nand NAND2_1273(g22845,g19441,g20885);
  nand NAND2_1274(g22846,g8278,g21660);
  nand NAND3_58(g22850,g21858,g21855,g21881);
  nand NAND2_1275(g22876,g21238,g83);
  nand NAND3_59(g22879,g21870,g21866,g21862);
  nand NAND2_1276(g22880,g19468,g20904);
  nand NAND2_1277(g22881,g8287,g21689);
  nand NAND3_60(g22885,g21863,g21859,g21885);
  nand NAND2_1278(g22911,g21246,g771);
  nand NAND3_61(g22914,g21874,g21871,g21868);
  nand NAND2_1279(g22915,g19491,g20928);
  nand NAND2_1280(g22916,g8296,g21725);
  nand NAND3_62(g22920,g21869,g21864,g21888);
  nand NAND2_1281(g22936,g21255,g1457);
  nand NAND3_63(g22939,g21877,g21875,g21873);
  nand NAND2_1282(g22940,g19512,g20956);
  nand NAND2_1283(g22941,g8305,g21751);
  nand NAND2_1284(g22942,g21263,g2151);
  nand NAND2_1285(g22992,g21636,g672);
  nand NAND2_1286(g23003,g21667,g1358);
  nand NAND2_1287(g23017,g21696,g2052);
  nand NAND2_1288(g23033,g21732,g2746);
  nand NAND2_1289(g23320,g23066,g23051);
  nand NAND2_1290(g23325,g23080,g23070);
  nand NAND2_1291(g23331,g22999,g22174);
  nand NAND2_1292(g23335,g23096,g23083);
  nand NAND2_1293(g23340,g23013,g22189);
  nand NAND2_1294(g23344,g23113,g23099);
  nand NAND2_1295(g23349,g23029,g22198);
  nand NAND2_1296(g23353,g23046,g22204);
  nand NAND2_1297(g23360,g21980,g21975);
  nand NAND2_1298(g23364,g21987,g21981);
  nand NAND2_1299(g23368,g23135,g22288);
  nand NAND2_1300(g23372,g22000,g21988);
  nand NAND2_1301(g23376,g18435,g22812);
  nand NAND2_1302(g23377,g21968,g22308);
  nand NAND2_1303(g23381,g22013,g22001);
  nand NAND2_1304(g23387,g18508,g22852);
  nand NAND2_1305(g23388,g21971,g22336);
  nand NAND2_1306(g23394,g18572,g22887);
  nand NAND2_1307(g23395,g21973,g22361);
  nand NAND2_1308(g23402,g18622,g22922);
  nand NAND3_64(g23478,g22809,g14442,g10694);
  nand NAND3_65(g23486,g22844,g14442,g10694);
  nand NAND3_66(g23489,g22850,g14529,g10714);
  nand NAND3_67(g23495,g10694,g14442,g22316);
  nand NAND3_68(g23502,g22879,g14529,g10714);
  nand NAND3_69(g23505,g22885,g14584,g10735);
  nand NAND3_70(g23511,g10714,g14529,g22341);
  nand NAND3_71(g23518,g22914,g14584,g10735);
  nand NAND3_72(g23521,g22920,g14618,g10754);
  nand NAND3_73(g23526,g10735,g14584,g22364);
  nand NAND3_74(g23533,g22939,g14618,g10754);
  nand NAND3_75(g23537,g10754,g14618,g22384);
  nand NAND2_1309(II30790,g22846,g14079);
  nand NAND2_1310(II30791,g22846,II30790);
  nand NAND2_1311(II30792,g14079,II30790);
  nand NAND2_1312(g23660,II30791,II30792);
  nand NAND2_1313(II30868,g22881,g14194);
  nand NAND2_1314(II30869,g22881,II30868);
  nand NAND2_1315(II30870,g14194,II30868);
  nand NAND2_1316(g23710,II30869,II30870);
  nand NAND2_1317(II30952,g22916,g14309);
  nand NAND2_1318(II30953,g22916,II30952);
  nand NAND2_1319(II30954,g14309,II30952);
  nand NAND2_1320(g23764,II30953,II30954);
  nand NAND2_1321(II31035,g22941,g14431);
  nand NAND2_1322(II31036,g22941,II31035);
  nand NAND2_1323(II31037,g14431,II31035);
  nand NAND2_1324(g23819,II31036,II31037);
  nand NAND2_1325(g23906,g22812,g13958);
  nand NAND2_1326(g23936,g22812,g13922);
  nand NAND2_1327(g23937,g22812,g13918);
  nand NAND2_1328(g23938,g22852,g14028);
  nand NAND2_1329(g23953,g22812,g14525);
  nand NAND2_1330(g23968,g22852,g13978);
  nand NAND2_1331(g23969,g22852,g13974);
  nand NAND2_1332(g23970,g22887,g14119);
  nand NAND2_1333(g23973,g22812,g14450);
  nand NAND2_1334(g23982,g22852,g14580);
  nand NAND2_1335(g23997,g22887,g14048);
  nand NAND2_1336(g23998,g22887,g14044);
  nand NAND2_1337(g23999,g22922,g14234);
  nand NAND2_1338(g24002,g22812,g14355);
  nand NAND2_1339(g24003,g22852,g14537);
  nand NAND2_1340(g24012,g22887,g14614);
  nand NAND2_1341(g24027,g22922,g14139);
  nand NAND2_1342(g24028,g22922,g14135);
  nand NAND2_1343(g24034,g22812,g14252);
  nand NAND2_1344(g24036,g22852,g14467);
  nand NAND2_1345(g24037,g22887,g14592);
  nand NAND2_1346(g24046,g22922,g14637);
  nand NAND2_1347(g24052,g22812,g14171);
  nand NAND2_1348(g24054,g22852,g14374);
  nand NAND2_1349(g24056,g22887,g14554);
  nand NAND2_1350(g24057,g22922,g14626);
  nand NAND2_1351(g24058,g22812,g14086);
  nand NAND2_1352(g24065,g22852,g14286);
  nand NAND2_1353(g24067,g22887,g14486);
  nand NAND2_1354(g24069,g22922,g14609);
  nand NAND2_1355(g24070,g22812,g14011);
  nand NAND2_1356(g24071,g22852,g14201);
  nand NAND2_1357(g24078,g22887,g14408);
  nand NAND2_1358(g24080,g22922,g14573);
  nand NAND2_1359(g24081,g22852,g14102);
  nand NAND2_1360(g24082,g22887,g14316);
  nand NAND2_1361(g24089,g22922,g14520);
  nand NAND2_1362(g24090,g22887,g14217);
  nand NAND2_1363(g24091,g22922,g14438);
  nand NAND2_1364(g24093,g22922,g14332);
  nand NAND2_1365(g24100,g20885,g22175);
  nand NAND2_1366(g24109,g20904,g22190);
  nand NAND2_1367(g24126,g20928,g22199);
  nand NAND2_1368(g24145,g20956,g22205);
  nand NAND2_1369(g24442,g23644,g3306);
  nand NAND2_1370(g24443,g23644,g3306);
  nand NAND2_1371(g24444,g23694,g3462);
  nand NAND2_1372(g24447,g23644,g3306);
  nand NAND2_1373(g24448,g23923,g3338);
  nand NAND2_1374(g24449,g23694,g3462);
  nand NAND2_1375(g24450,g23748,g3618);
  nand NAND2_1376(g24451,g23644,g3306);
  nand NAND2_1377(g24452,g23923,g3338);
  nand NAND2_1378(g24453,g23694,g3462);
  nand NAND2_1379(g24454,g23955,g3494);
  nand NAND2_1380(g24455,g23748,g3618);
  nand NAND2_1381(g24456,g23803,g3774);
  nand NAND2_1382(g24457,g23923,g3338);
  nand NAND2_1383(g24458,g23694,g3462);
  nand NAND2_1384(g24459,g23955,g3494);
  nand NAND2_1385(g24460,g23748,g3618);
  nand NAND2_1386(g24461,g23984,g3650);
  nand NAND2_1387(g24462,g23803,g3774);
  nand NAND2_1388(g24463,g23923,g3338);
  nand NAND2_1389(g24464,g23955,g3494);
  nand NAND2_1390(g24465,g23748,g3618);
  nand NAND2_1391(g24466,g23984,g3650);
  nand NAND2_1392(g24467,g23803,g3774);
  nand NAND2_1393(g24468,g24014,g3806);
  nand NAND2_1394(g24469,g23955,g3494);
  nand NAND2_1395(g24470,g23984,g3650);
  nand NAND2_1396(g24471,g23803,g3774);
  nand NAND2_1397(g24472,g24014,g3806);
  nand NAND2_1398(g24474,g23984,g3650);
  nand NAND2_1399(g24475,g24014,g3806);
  nand NAND2_1400(g24477,g24014,g3806);
  nand NAND2_1401(g24616,g499,g23376);
  nand NAND2_1402(g24627,g1186,g23387);
  nand NAND2_1403(g24641,g1880,g23394);
  nand NAND2_1404(g24660,g2574,g23402);
  nand NAND2_1405(II32265,g17903,g23936);
  nand NAND2_1406(II32266,g17903,II32265);
  nand NAND2_1407(II32267,g23936,II32265);
  nand NAND2_1408(g24753,II32266,II32267);
  nand NAND2_1409(II32284,g17815,g23953);
  nand NAND2_1410(II32285,g17815,II32284);
  nand NAND2_1411(II32286,g23953,II32284);
  nand NAND2_1412(g24766,II32285,II32286);
  nand NAND2_1413(II32295,g18014,g23968);
  nand NAND2_1414(II32296,g18014,II32295);
  nand NAND2_1415(II32297,g23968,II32295);
  nand NAND2_1416(g24771,II32296,II32297);
  nand NAND2_1417(II32308,g17903,g23973);
  nand NAND2_1418(II32309,g17903,II32308);
  nand NAND2_1419(II32310,g23973,II32308);
  nand NAND2_1420(g24778,II32309,II32310);
  nand NAND2_1421(II32323,g17927,g23982);
  nand NAND2_1422(II32324,g17927,II32323);
  nand NAND2_1423(II32325,g23982,II32323);
  nand NAND2_1424(g24787,II32324,II32325);
  nand NAND2_1425(II32333,g18131,g23997);
  nand NAND2_1426(II32334,g18131,II32333);
  nand NAND2_1427(II32335,g23997,II32333);
  nand NAND2_1428(g24791,II32334,II32335);
  nand NAND2_1429(II32345,g17815,g24002);
  nand NAND2_1430(II32346,g17815,II32345);
  nand NAND2_1431(II32347,g24002,II32345);
  nand NAND2_1432(g24797,II32346,II32347);
  nand NAND2_1433(II32355,g18014,g24003);
  nand NAND2_1434(II32356,g18014,II32355);
  nand NAND2_1435(II32357,g24003,II32355);
  nand NAND2_1436(g24801,II32356,II32357);
  nand NAND2_1437(II32368,g18038,g24012);
  nand NAND2_1438(II32369,g18038,II32368);
  nand NAND2_1439(II32370,g24012,II32368);
  nand NAND2_1440(g24808,II32369,II32370);
  nand NAND2_1441(II32378,g18247,g24027);
  nand NAND2_1442(II32379,g18247,II32378);
  nand NAND2_1443(II32380,g24027,II32378);
  nand NAND2_1444(g24812,II32379,II32380);
  nand NAND2_1445(g24814,g24239,g24244);
  nand NAND2_1446(II32391,g17903,g24034);
  nand NAND2_1447(II32392,g17903,II32391);
  nand NAND2_1448(II32393,g24034,II32391);
  nand NAND2_1449(g24817,II32392,II32393);
  nand NAND2_1450(II32400,g17927,g24036);
  nand NAND2_1451(II32401,g17927,II32400);
  nand NAND2_1452(II32402,g24036,II32400);
  nand NAND2_1453(g24820,II32401,II32402);
  nand NAND2_1454(II32409,g18131,g24037);
  nand NAND2_1455(II32410,g18131,II32409);
  nand NAND2_1456(II32411,g24037,II32409);
  nand NAND2_1457(g24823,II32410,II32411);
  nand NAND2_1458(II32422,g18155,g24046);
  nand NAND2_1459(II32423,g18155,II32422);
  nand NAND2_1460(II32424,g24046,II32422);
  nand NAND2_1461(g24830,II32423,II32424);
  nand NAND2_1462(II32430,g17815,g24052);
  nand NAND2_1463(II32431,g17815,II32430);
  nand NAND2_1464(II32432,g24052,II32430);
  nand NAND2_1465(g24832,II32431,II32432);
  nand NAND2_1466(g24833,g24245,g24252);
  nand NAND2_1467(II32443,g18014,g24054);
  nand NAND2_1468(II32444,g18014,II32443);
  nand NAND2_1469(II32445,g24054,II32443);
  nand NAND2_1470(g24837,II32444,II32445);
  nand NAND2_1471(II32451,g18038,g24056);
  nand NAND2_1472(II32452,g18038,II32451);
  nand NAND2_1473(II32453,g24056,II32451);
  nand NAND2_1474(g24839,II32452,II32453);
  nand NAND2_1475(II32460,g18247,g24057);
  nand NAND2_1476(II32461,g18247,II32460);
  nand NAND2_1477(II32462,g24057,II32460);
  nand NAND2_1478(g24842,II32461,II32462);
  nand NAND2_1479(II32468,g17903,g24058);
  nand NAND2_1480(II32469,g17903,II32468);
  nand NAND2_1481(II32470,g24058,II32468);
  nand NAND2_1482(g24844,II32469,II32470);
  nand NAND2_1483(II32478,g17927,g24065);
  nand NAND2_1484(II32479,g17927,II32478);
  nand NAND2_1485(II32480,g24065,II32478);
  nand NAND2_1486(g24848,II32479,II32480);
  nand NAND2_1487(g24849,g24254,g24257);
  nand NAND2_1488(II32490,g18131,g24067);
  nand NAND2_1489(II32491,g18131,II32490);
  nand NAND2_1490(II32492,g24067,II32490);
  nand NAND2_1491(g24852,II32491,II32492);
  nand NAND2_1492(II32498,g18155,g24069);
  nand NAND2_1493(II32499,g18155,II32498);
  nand NAND2_1494(II32500,g24069,II32498);
  nand NAND2_1495(g24854,II32499,II32500);
  nand NAND2_1496(II32509,g17815,g24070);
  nand NAND2_1497(II32510,g17815,II32509);
  nand NAND2_1498(II32511,g24070,II32509);
  nand NAND2_1499(g24857,II32510,II32511);
  nand NAND2_1500(II32518,g18014,g24071);
  nand NAND2_1501(II32519,g18014,II32518);
  nand NAND2_1502(II32520,g24071,II32518);
  nand NAND2_1503(g24860,II32519,II32520);
  nand NAND2_1504(II32526,g18038,g24078);
  nand NAND2_1505(II32527,g18038,II32526);
  nand NAND2_1506(II32528,g24078,II32526);
  nand NAND2_1507(g24862,II32527,II32528);
  nand NAND2_1508(g24863,g24258,g23319);
  nand NAND2_1509(II32538,g18247,g24080);
  nand NAND2_1510(II32539,g18247,II32538);
  nand NAND2_1511(II32540,g24080,II32538);
  nand NAND2_1512(g24866,II32539,II32540);
  nand NAND2_1513(II32546,g17903,g23906);
  nand NAND2_1514(II32547,g17903,II32546);
  nand NAND2_1515(II32548,g23906,II32546);
  nand NAND2_1516(g24868,II32547,II32548);
  nand NAND2_1517(II32559,g17927,g24081);
  nand NAND2_1518(II32560,g17927,II32559);
  nand NAND2_1519(II32561,g24081,II32559);
  nand NAND2_1520(g24873,II32560,II32561);
  nand NAND2_1521(II32567,g18131,g24082);
  nand NAND2_1522(II32568,g18131,II32567);
  nand NAND2_1523(II32569,g24082,II32567);
  nand NAND2_1524(g24875,II32568,II32569);
  nand NAND2_1525(II32575,g18155,g24089);
  nand NAND2_1526(II32576,g18155,II32575);
  nand NAND2_1527(II32577,g24089,II32575);
  nand NAND2_1528(g24877,II32576,II32577);
  nand NAND2_1529(II32586,g17815,g23937);
  nand NAND2_1530(II32587,g17815,II32586);
  nand NAND2_1531(II32588,g23937,II32586);
  nand NAND2_1532(g24880,II32587,II32588);
  nand NAND2_1533(II32595,g18014,g23938);
  nand NAND2_1534(II32596,g18014,II32595);
  nand NAND2_1535(II32597,g23938,II32595);
  nand NAND2_1536(g24883,II32596,II32597);
  nand NAND2_1537(II32607,g18038,g24090);
  nand NAND2_1538(II32608,g18038,II32607);
  nand NAND2_1539(II32609,g24090,II32607);
  nand NAND2_1540(g24887,II32608,II32609);
  nand NAND2_1541(II32615,g18247,g24091);
  nand NAND2_1542(II32616,g18247,II32615);
  nand NAND2_1543(II32617,g24091,II32615);
  nand NAND2_1544(g24889,II32616,II32617);
  nand NAND2_1545(II32624,g17927,g23969);
  nand NAND2_1546(II32625,g17927,II32624);
  nand NAND2_1547(II32626,g23969,II32624);
  nand NAND2_1548(g24897,II32625,II32626);
  nand NAND2_1549(II32633,g18131,g23970);
  nand NAND2_1550(II32634,g18131,II32633);
  nand NAND2_1551(II32635,g23970,II32633);
  nand NAND2_1552(g24900,II32634,II32635);
  nand NAND2_1553(II32645,g18155,g24093);
  nand NAND2_1554(II32646,g18155,II32645);
  nand NAND2_1555(II32647,g24093,II32645);
  nand NAND2_1556(g24904,II32646,II32647);
  nand NAND2_1557(II32659,g18038,g23998);
  nand NAND2_1558(II32660,g18038,II32659);
  nand NAND2_1559(II32661,g23998,II32659);
  nand NAND2_1560(g24920,II32660,II32661);
  nand NAND2_1561(II32668,g18247,g23999);
  nand NAND2_1562(II32669,g18247,II32668);
  nand NAND2_1563(II32670,g23999,II32668);
  nand NAND2_1564(g24923,II32669,II32670);
  nand NAND2_1565(II32677,g23823,g14165);
  nand NAND2_1566(II32678,g23823,II32677);
  nand NAND2_1567(II32679,g14165,II32677);
  nand NAND2_1568(g24928,II32678,II32679);
  nand NAND2_1569(II32686,g18155,g24028);
  nand NAND2_1570(II32687,g18155,II32686);
  nand NAND2_1571(II32688,g24028,II32686);
  nand NAND2_1572(g24937,II32687,II32688);
  nand NAND2_1573(II32695,g23858,g14280);
  nand NAND2_1574(II32696,g23858,II32695);
  nand NAND2_1575(II32697,g14280,II32695);
  nand NAND2_1576(g24940,II32696,II32697);
  nand NAND2_1577(II32708,g23892,g14402);
  nand NAND2_1578(II32709,g23892,II32708);
  nand NAND2_1579(II32710,g14402,II32708);
  nand NAND2_1580(g24951,II32709,II32710);
  nand NAND2_1581(II32724,g23913,g14514);
  nand NAND2_1582(II32725,g23913,II32724);
  nand NAND2_1583(II32726,g14514,II32724);
  nand NAND2_1584(g24963,II32725,II32726);
  nand NAND2_1585(g24975,g23497,g74);
  nand NAND2_1586(g24986,g23513,g762);
  nand NAND2_1587(g24997,g23528,g1448);
  nand NAND2_1588(g25004,g23644,g6448);
  nand NAND2_1589(g25005,g23539,g2142);
  nand NAND2_1590(g25008,g23644,g5438);
  nand NAND2_1591(g25009,g23644,g6448);
  nand NAND2_1592(g25010,g23694,g6713);
  nand NAND2_1593(g25011,g23644,g5438);
  nand NAND2_1594(g25012,g23644,g6448);
  nand NAND2_1595(g25013,g23923,g6643);
  nand NAND2_1596(g25014,g23694,g5473);
  nand NAND2_1597(g25015,g23694,g6713);
  nand NAND2_1598(g25016,g23748,g7015);
  nand NAND2_1599(g25017,g23644,g5438);
  nand NAND2_1600(g25018,g23644,g6448);
  nand NAND2_1601(g25019,g23923,g6486);
  nand NAND2_1602(g25020,g23923,g6643);
  nand NAND2_1603(g25021,g23694,g5473);
  nand NAND2_1604(g25022,g23694,g6713);
  nand NAND2_1605(g25023,g23955,g6945);
  nand NAND2_1606(g25024,g23748,g5512);
  nand NAND2_1607(g25025,g23748,g7015);
  nand NAND2_1608(g25026,g23803,g7265);
  nand NAND2_1609(g25028,g23644,g5438);
  nand NAND2_1610(g25029,g23923,g6486);
  nand NAND2_1611(g25030,g23923,g6643);
  nand NAND2_1612(g25031,g23694,g5473);
  nand NAND2_1613(g25032,g23694,g6713);
  nand NAND2_1614(g25033,g23955,g6751);
  nand NAND2_1615(g25034,g23955,g6945);
  nand NAND2_1616(g25035,g23748,g5512);
  nand NAND2_1617(g25036,g23748,g7015);
  nand NAND2_1618(g25037,g23984,g7195);
  nand NAND2_1619(g25038,g23803,g5556);
  nand NAND2_1620(g25039,g23803,g7265);
  nand NAND2_1621(g25040,g23923,g6486);
  nand NAND2_1622(g25041,g23923,g6643);
  nand NAND2_1623(g25043,g23694,g5473);
  nand NAND2_1624(g25044,g23955,g6751);
  nand NAND2_1625(g25045,g23955,g6945);
  nand NAND2_1626(g25046,g23748,g5512);
  nand NAND2_1627(g25047,g23748,g7015);
  nand NAND2_1628(g25048,g23984,g7053);
  nand NAND2_1629(g25049,g23984,g7195);
  nand NAND2_1630(g25050,g23803,g5556);
  nand NAND2_1631(g25051,g23803,g7265);
  nand NAND2_1632(g25052,g24014,g7391);
  nand NAND2_1633(g25053,g23923,g6486);
  nand NAND2_1634(g25054,g23955,g6751);
  nand NAND2_1635(g25055,g23955,g6945);
  nand NAND2_1636(g25057,g23748,g5512);
  nand NAND2_1637(g25058,g23984,g7053);
  nand NAND2_1638(g25059,g23984,g7195);
  nand NAND2_1639(g25060,g23803,g5556);
  nand NAND2_1640(g25061,g23803,g7265);
  nand NAND2_1641(g25062,g24014,g7303);
  nand NAND2_1642(g25063,g24014,g7391);
  nand NAND2_1643(g25064,g23955,g6751);
  nand NAND2_1644(g25065,g23984,g7053);
  nand NAND2_1645(g25066,g23984,g7195);
  nand NAND2_1646(g25068,g23803,g5556);
  nand NAND2_1647(g25069,g24014,g7303);
  nand NAND2_1648(g25070,g24014,g7391);
  nand NAND2_1649(g25071,g23984,g7053);
  nand NAND2_1650(g25072,g24014,g7303);
  nand NAND2_1651(g25073,g24014,g7391);
  nand NAND2_1652(g25074,g24014,g7303);
  nand NAND2_1653(g25088,g23950,g679);
  nand NAND2_1654(g25096,g23979,g1365);
  nand NAND2_1655(g25106,g24009,g2059);
  nand NAND2_1656(g25112,g24043,g2753);
  nand NAND2_1657(g25200,g24965,g3306);
  nand NAND2_1658(g25203,g24978,g3462);
  nand NAND2_1659(g25205,g24989,g3618);
  nand NAND2_1660(g25210,g25000,g3774);
  nand NAND4_5(g25312,g21211,g14442,g10694,g24590);
  nand NAND4_6(g25320,g21219,g14529,g10714,g24595);
  nand NAND4_7(g25331,g21230,g14584,g10735,g24603);
  nand NAND4_8(g25340,g21235,g14618,g10754,g24610);
  nand NAND2_1661(g25927,g24965,g6448);
  nand NAND2_1662(g25928,g24965,g5438);
  nand NAND2_1663(g25929,g24978,g6713);
  nand NAND2_1664(g25930,g24978,g5473);
  nand NAND2_1665(g25931,g24989,g7015);
  nand NAND2_1666(g25933,g24989,g5512);
  nand NAND2_1667(g25934,g25000,g7265);
  nand NAND2_1668(g25936,g25000,g5556);
  nand NAND2_1669(g25954,g22806,g24517);
  nand NAND2_1670(g25958,g22847,g24530);
  nand NAND2_1671(g25964,g22882,g24543);
  nand NAND2_1672(g25969,g22917,g24555);
  nand NAND3_76(g26059,g25422,g25379,g25274);
  nand NAND3_77(g26066,g25431,g25395,g25283);
  nand NAND3_78(g26073,g25438,g25405,g25291);
  nand NAND3_79(g26079,g25445,g25413,g25301);
  nand NAND2_1673(g26106,g23644,g25354);
  nand NAND4_9(g26119,g8278,g14657,g25422,g25379);
  nand NAND2_1674(g26120,g23694,g25369);
  nand NAND4_10(g26129,g8287,g14691,g25431,g25395);
  nand NAND2_1675(g26130,g23748,g25386);
  nand NAND4_11(g26143,g8296,g14725,g25438,g25405);
  nand NAND2_1676(g26144,g23803,g25402);
  nand NAND4_12(g26148,g8305,g14753,g25445,g25413);
  nand NAND2_1677(g26356,g16539,g25183);
  nand NAND2_1678(g26399,g16571,g25186);
  nand NAND2_1679(g26440,g16595,g25190);
  nand NAND2_1680(g26458,g25343,g65);
  nand NAND2_1681(g26472,g16615,g25195);
  nand NAND2_1682(g26482,g25357,g753);
  nand NAND2_1683(g26498,g25372,g1439);
  nand NAND2_1684(g26513,g25389,g2133);
  nand NAND2_1685(g26772,g26320,g3306);
  nand NAND2_1686(g26779,g26367,g3462);
  nand NAND2_1687(g26785,g26410,g3618);
  nand NAND2_1688(g26792,g26451,g3774);
  nand NAND2_1689(II35020,g26110,g26099);
  nand NAND2_1690(II35021,g26110,II35020);
  nand NAND2_1691(II35022,g26099,II35020);
  nand NAND2_1692(g26859,II35021,II35022);
  nand NAND2_1693(II35034,g26087,g26154);
  nand NAND2_1694(II35035,g26087,II35034);
  nand NAND2_1695(II35036,g26154,II35034);
  nand NAND2_1696(g26865,II35035,II35036);
  nand NAND2_1697(II35042,g26151,g26145);
  nand NAND2_1698(II35043,g26151,II35042);
  nand NAND2_1699(II35044,g26145,II35042);
  nand NAND2_1700(g26867,II35043,II35044);
  nand NAND2_1701(II35057,g26137,g26126);
  nand NAND2_1702(II35058,g26137,II35057);
  nand NAND2_1703(II35059,g26126,II35057);
  nand NAND2_1704(g26874,II35058,II35059);
  nand NAND4_13(g26892,g25699,g26283,g25569,g25631);
  nand NAND3_80(g26902,g25631,g26283,g25569);
  nand NAND4_14(g26906,g25772,g26327,g25648,g25708);
  nand NAND2_1705(g26911,g25569,g26283);
  nand NAND3_81(g26915,g25708,g26327,g25648);
  nand NAND4_15(g26918,g25826,g26374,g25725,g25781);
  nand NAND2_1706(g26925,g25648,g26327);
  nand NAND3_82(g26928,g25781,g26374,g25725);
  nand NAND4_16(g26931,g25861,g26417,g25798,g25835);
  nand NAND2_1707(II35123,g26107,g26096);
  nand NAND2_1708(II35124,g26107,II35123);
  nand NAND2_1709(II35125,g26096,II35123);
  nand NAND2_1710(g26934,II35124,II35125);
  nand NAND2_1711(g26938,g25725,g26374);
  nand NAND3_83(g26941,g25835,g26417,g25798);
  nand NAND2_1712(g26947,g25798,g26417);
  nand NAND2_1713(g27117,g26320,g6448);
  nand NAND2_1714(g27118,g26320,g5438);
  nand NAND2_1715(g27119,g26367,g6713);
  nand NAND2_1716(g27121,g26367,g5473);
  nand NAND2_1717(g27122,g26410,g7015);
  nand NAND2_1718(g27124,g26410,g5512);
  nand NAND2_1719(g27125,g26451,g7265);
  nand NAND2_1720(g27130,g26451,g5556);
  nand NAND2_1721(II35701,g26867,g26874);
  nand NAND2_1722(II35702,g26867,II35701);
  nand NAND2_1723(II35703,g26874,II35701);
  nand NAND2_1724(g27379,II35702,II35703);
  nand NAND2_1725(II35714,g26859,g26865);
  nand NAND2_1726(II35715,g26859,II35714);
  nand NAND2_1727(II35716,g26865,II35714);
  nand NAND2_1728(g27382,II35715,II35716);
  nand NAND2_1729(g27390,g26989,g6448);
  nand NAND2_1730(g27395,g26989,g5438);
  nand NAND2_1731(g27400,g27012,g6713);
  nand NAND2_1732(g27408,g27012,g5473);
  nand NAND2_1733(g27413,g27038,g7015);
  nand NAND2_1734(g27426,g27038,g5512);
  nand NAND2_1735(g27431,g27066,g7265);
  nand NAND2_1736(g27447,g27066,g5556);
  nand NAND2_1737(II35904,g27051,g14831);
  nand NAND2_1738(II35905,g27051,II35904);
  nand NAND2_1739(II35906,g14831,II35904);
  nand NAND2_1740(g27528,II35905,II35906);
  nand NAND2_1741(II35944,g27078,g14904);
  nand NAND2_1742(II35945,g27078,II35944);
  nand NAND2_1743(II35946,g14904,II35944);
  nand NAND2_1744(g27550,II35945,II35946);
  nand NAND2_1745(II35974,g27094,g14985);
  nand NAND2_1746(II35975,g27094,II35974);
  nand NAND2_1747(II35976,g14985,II35974);
  nand NAND2_1748(g27566,II35975,II35976);
  nand NAND2_1749(g27571,g26869,g56);
  nand NAND2_1750(II35992,g27106,g15074);
  nand NAND2_1751(II35993,g27106,II35992);
  nand NAND2_1752(II35994,g15074,II35992);
  nand NAND2_1753(g27576,II35993,II35994);
  nand NAND2_1754(g27580,g26878,g744);
  nand NAND2_1755(g27583,g26887,g1430);
  nand NAND2_1756(g27587,g26897,g2124);
  nand NAND2_1757(g27626,g26989,g3306);
  nand NAND2_1758(g27627,g27012,g3462);
  nand NAND2_1759(g27628,g27038,g3618);
  nand NAND2_1760(g27630,g27066,g3774);
  nand NAND2_1761(g27738,g25367,g27415);
  nand NAND2_1762(g27743,g25384,g27436);
  nand NAND2_1763(g27751,g25400,g27455);
  nand NAND2_1764(g27756,g25410,g27471);
  nand NAND2_1765(II36256,g27527,g15859);
  nand NAND2_1766(II36257,g27527,II36256);
  nand NAND2_1767(II36258,g15859,II36256);
  nand NAND2_1768(g27801,II36257,II36258);
  nand NAND2_1769(II36270,g27549,g15890);
  nand NAND2_1770(II36271,g27549,II36270);
  nand NAND2_1771(II36272,g15890,II36270);
  nand NAND2_1772(g27809,II36271,II36272);
  nand NAND2_1773(II36289,g27565,g15923);
  nand NAND2_1774(II36290,g27565,II36289);
  nand NAND2_1775(II36291,g15923,II36289);
  nand NAND2_1776(g27830,II36290,II36291);
  nand NAND2_1777(II36300,g27382,g27379);
  nand NAND2_1778(II36301,g27382,II36300);
  nand NAND2_1779(II36302,g27379,II36300);
  nand NAND2_1780(g27838,II36301,II36302);
  nand NAND2_1781(II36314,g27575,g15952);
  nand NAND2_1782(II36315,g27575,II36314);
  nand NAND2_1783(II36316,g15952,II36314);
  nand NAND2_1784(g27846,II36315,II36316);
  nand NAND2_1785(II36591,g27529,g14885);
  nand NAND2_1786(II36592,g27529,II36591);
  nand NAND2_1787(II36593,g14885,II36591);
  nand NAND2_1788(g28046,II36592,II36593);
  nand NAND2_1789(II36666,g27551,g14966);
  nand NAND2_1790(II36667,g27551,II36666);
  nand NAND2_1791(II36668,g14966,II36666);
  nand NAND2_1792(g28075,II36667,II36668);
  nand NAND2_1793(II36731,g27567,g15055);
  nand NAND2_1794(II36732,g27567,II36731);
  nand NAND2_1795(II36733,g15055,II36731);
  nand NAND2_1796(g28100,II36732,II36733);
  nand NAND2_1797(II36779,g27577,g15151);
  nand NAND2_1798(II36780,g27577,II36779);
  nand NAND2_1799(II36781,g15151,II36779);
  nand NAND2_1800(g28118,II36780,II36781);
  nand NAND2_1801(II37295,g27827,g27814);
  nand NAND2_1802(II37296,g27827,II37295);
  nand NAND2_1803(II37297,g27814,II37295);
  nand NAND2_1804(g28384,II37296,II37297);
  nand NAND2_1805(II37303,g27802,g27900);
  nand NAND2_1806(II37304,g27802,II37303);
  nand NAND2_1807(II37305,g27900,II37303);
  nand NAND2_1808(g28386,II37304,II37305);
  nand NAND2_1809(II37311,g27897,g27883);
  nand NAND2_1810(II37312,g27897,II37311);
  nand NAND2_1811(II37313,g27883,II37311);
  nand NAND2_1812(g28388,II37312,II37313);
  nand NAND2_1813(II37322,g27865,g27855);
  nand NAND2_1814(II37323,g27865,II37322);
  nand NAND2_1815(II37324,g27855,II37322);
  nand NAND2_1816(g28391,II37323,II37324);
  nand NAND2_1817(II37356,g27824,g27811);
  nand NAND2_1818(II37357,g27824,II37356);
  nand NAND2_1819(II37358,g27811,II37356);
  nand NAND2_1820(g28415,II37357,II37358);
  nand NAND2_1821(II37813,g28388,g28391);
  nand NAND2_1822(II37814,g28388,II37813);
  nand NAND2_1823(II37815,g28391,II37813);
  nand NAND2_1824(g28842,II37814,II37815);
  nand NAND2_1825(II37822,g28384,g28386);
  nand NAND2_1826(II37823,g28384,II37822);
  nand NAND2_1827(II37824,g28386,II37822);
  nand NAND2_1828(g28845,II37823,II37824);
  nand NAND2_1829(g28978,g9150,g28512);
  nand NAND2_1830(g29001,g9161,g28512);
  nand NAND2_1831(g29008,g9174,g28540);
  nand NAND2_1832(g29026,g9187,g28512);
  nand NAND2_1833(g29030,g9203,g28540);
  nand NAND2_1834(g29038,g9216,g28567);
  nand NAND2_1835(g29045,g9232,g28512);
  nand NAND2_1836(g29049,g9248,g28540);
  nand NAND2_1837(g29053,g9264,g28567);
  nand NAND2_1838(g29060,g9277,g28595);
  nand NAND2_1839(g29062,g9310,g28540);
  nand NAND2_1840(g29068,g9326,g28567);
  nand NAND2_1841(g29072,g9342,g28595);
  nand NAND2_1842(g29076,g9391,g28567);
  nand NAND2_1843(g29080,g9407,g28595);
  nand NAND2_1844(g29087,g9488,g28595);
  nand NAND2_1845(g29088,g9507,g28512);
  nand NAND2_1846(g29096,g9649,g28540);
  nand NAND2_1847(g29103,g9795,g28567);
  nand NAND2_1848(g29107,g9941,g28595);
  nand NAND2_1849(II38378,g28845,g28842);
  nand NAND2_1850(II38379,g28845,II38378);
  nand NAND2_1851(II38380,g28842,II38378);
  nand NAND2_1852(g29265,II38379,II38380);
  nand NAND2_1853(II38810,g29303,g15904);
  nand NAND2_1854(II38811,g29303,II38810);
  nand NAND2_1855(II38812,g15904,II38810);
  nand NAND2_1856(g29498,II38811,II38812);
  nand NAND2_1857(II38820,g29313,g15933);
  nand NAND2_1858(II38821,g29313,II38820);
  nand NAND2_1859(II38822,g15933,II38820);
  nand NAND2_1860(g29500,II38821,II38822);
  nand NAND2_1861(II38831,g29324,g15962);
  nand NAND2_1862(II38832,g29324,II38831);
  nand NAND2_1863(II38833,g15962,II38831);
  nand NAND2_1864(g29503,II38832,II38833);
  nand NAND2_1865(II38841,g29333,g15981);
  nand NAND2_1866(II38842,g29333,II38841);
  nand NAND2_1867(II38843,g15981,II38841);
  nand NAND2_1868(g29505,II38842,II38843);
  nand NAND2_1869(II39323,g29721,g29713);
  nand NAND2_1870(II39324,g29721,II39323);
  nand NAND2_1871(II39325,g29713,II39323);
  nand NAND2_1872(g29911,II39324,II39325);
  nand NAND2_1873(II39331,g29705,g29751);
  nand NAND2_1874(II39332,g29705,II39331);
  nand NAND2_1875(II39333,g29751,II39331);
  nand NAND2_1876(g29913,II39332,II39333);
  nand NAND2_1877(II39339,g29748,g29741);
  nand NAND2_1878(II39340,g29748,II39339);
  nand NAND2_1879(II39341,g29741,II39339);
  nand NAND2_1880(g29915,II39340,II39341);
  nand NAND2_1881(II39347,g29732,g29728);
  nand NAND2_1882(II39348,g29732,II39347);
  nand NAND2_1883(II39349,g29728,II39347);
  nand NAND2_1884(g29917,II39348,II39349);
  nand NAND2_1885(II39359,g29766,g15880);
  nand NAND2_1886(II39360,g29766,II39359);
  nand NAND2_1887(II39361,g15880,II39359);
  nand NAND2_1888(g29923,II39360,II39361);
  nand NAND2_1889(II39367,g29767,g15913);
  nand NAND2_1890(II39368,g29767,II39367);
  nand NAND2_1891(II39369,g15913,II39367);
  nand NAND2_1892(g29925,II39368,II39369);
  nand NAND2_1893(II39375,g29768,g15942);
  nand NAND2_1894(II39376,g29768,II39375);
  nand NAND2_1895(II39377,g15942,II39375);
  nand NAND2_1896(g29927,II39376,II39377);
  nand NAND2_1897(II39384,g29718,g29710);
  nand NAND2_1898(II39385,g29718,II39384);
  nand NAND2_1899(II39386,g29710,II39384);
  nand NAND2_1900(g29930,II39385,II39386);
  nand NAND2_1901(II39391,g29769,g15971);
  nand NAND2_1902(II39392,g29769,II39391);
  nand NAND2_1903(II39393,g15971,II39391);
  nand NAND2_1904(g29931,II39392,II39393);
  nand NAND2_1905(II39532,g29915,g29917);
  nand NAND2_1906(II39533,g29915,II39532);
  nand NAND2_1907(II39534,g29917,II39532);
  nand NAND2_1908(g30034,II39533,II39534);
  nand NAND2_1909(II39539,g29911,g29913);
  nand NAND2_1910(II39540,g29911,II39539);
  nand NAND2_1911(II39541,g29913,II39539);
  nand NAND2_1912(g30035,II39540,II39541);
  nand NAND2_1913(II39689,g30035,g30034);
  nand NAND2_1914(II39690,g30035,II39689);
  nand NAND2_1915(II39691,g30034,II39689);
  nand NAND2_1916(g30228,II39690,II39691);
  nand NAND2_1917(II40558,g30605,g30597);
  nand NAND2_1918(II40559,g30605,II40558);
  nand NAND2_1919(II40560,g30597,II40558);
  nand NAND2_1920(g30768,II40559,II40560);
  nand NAND2_1921(II40571,g30588,g30632);
  nand NAND2_1922(II40572,g30588,II40571);
  nand NAND2_1923(II40573,g30632,II40571);
  nand NAND2_1924(g30771,II40572,II40573);
  nand NAND2_1925(II40587,g30629,g30622);
  nand NAND2_1926(II40588,g30629,II40587);
  nand NAND2_1927(II40589,g30622,II40587);
  nand NAND2_1928(g30775,II40588,II40589);
  nand NAND2_1929(II40603,g30614,g30610);
  nand NAND2_1930(II40604,g30614,II40603);
  nand NAND2_1931(II40605,g30610,II40603);
  nand NAND2_1932(g30779,II40604,II40605);
  nand NAND2_1933(II40627,g30602,g30594);
  nand NAND2_1934(II40628,g30602,II40627);
  nand NAND2_1935(II40629,g30594,II40627);
  nand NAND2_1936(g30791,II40628,II40629);
  nand NAND2_1937(II41010,g30775,g30779);
  nand NAND2_1938(II41011,g30775,II41010);
  nand NAND2_1939(II41012,g30779,II41010);
  nand NAND2_1940(g30926,II41011,II41012);
  nand NAND2_1941(II41017,g30768,g30771);
  nand NAND2_1942(II41018,g30768,II41017);
  nand NAND2_1943(II41019,g30771,II41017);
  nand NAND2_1944(g30927,II41018,II41019);
  nand NAND2_1945(II41064,g30927,g30926);
  nand NAND2_1946(II41065,g30927,II41064);
  nand NAND2_1947(II41066,g30926,II41064);
  nand NAND2_1948(g30952,II41065,II41066);
  nor NOR3_0(g7528,g3151,g3142,g3147);
  nor NOR2_0(g7575,g2984,g2985);
  nor NOR2_1(g7795,g2992,g2991);
  nor NOR4_0(g8430,g3198,g8120,g3194,g3191);
  nor NOR3_1(g10784,g5630,g5649,g5676);
  nor NOR3_2(g10789,g5650,g5677,g5709);
  nor NOR3_3(g10793,g5658,g5687,g5728);
  nor NOR3_4(g10797,g5678,g5710,g5757);
  nor NOR3_5(g10801,g5688,g5729,g5767);
  nor NOR3_6(g10805,g5696,g5739,g5786);
  nor NOR3_7(g10810,g5711,g5758,g5807);
  nor NOR3_8(g10814,g5730,g5768,g5816);
  nor NOR3_9(g10818,g5740,g5787,g5826);
  nor NOR3_10(g10822,g5748,g5797,g5845);
  nor NOR3_11(g10831,g5769,g5817,g5863);
  nor NOR3_12(g10835,g5788,g5827,g5872);
  nor NOR3_13(g10839,g5798,g5846,g5882);
  nor NOR3_14(g10851,g5828,g5873,g5910);
  nor NOR3_15(g10855,g5847,g5883,g5919);
  nor NOR3_16(g10872,g5884,g5920,g5949);
  nor NOR3_17(g11600,g9049,g9064,g9078);
  nor NOR4_1(g11622,g8183,g11332,g7928,g11069);
  nor NOR3_18(g11624,g9062,g9075,g9091);
  nor NOR3_19(g11627,g9063,g9077,g9093);
  nor NOR3_20(g11630,g9066,g9081,g9097);
  nor NOR4_2(g11643,g11481,g8045,g7928,g11069);
  nor NOR3_21(g11644,g9076,g9092,g9102);
  nor NOR3_22(g11647,g9079,g9094,g9103);
  nor NOR3_23(g11650,g9080,g9096,g9105);
  nor NOR3_24(g11653,g9083,g9100,g9109);
  nor NOR4_3(g11660,g8183,g8045,g7928,g11069);
  nor NOR3_25(g11663,g9095,g9104,g9112);
  nor NOR3_26(g11666,g9098,g9106,g9113);
  nor NOR3_27(g11669,g9099,g9108,g9115);
  nor NOR3_28(g11675,g9107,g9114,g9120);
  nor NOR3_29(g11678,g9110,g9116,g9121);
  nor NOR3_30(g11681,g9111,g9118,g9123);
  nor NOR3_31(g11687,g9117,g9122,g9126);
  nor NOR3_32(g11690,g9119,g9124,g9127);
  nor NOR3_33(g11697,g9125,g9131,g9133);
  nor NOR3_34(g11703,g9132,g9137,g9139);
  nor NOR3_35(g11711,g9138,g9143,g9145);
  nor NOR3_36(g11744,g9241,g9301,g9364);
  nor NOR3_37(g11759,g9302,g9365,g9438);
  nor NOR3_38(g11760,g9319,g9382,g9461);
  nor NOR3_39(g11767,g9366,g9439,g9518);
  nor NOR3_40(g11768,g9367,g9441,g9521);
  nor NOR3_41(g11772,g9383,g9462,g9580);
  nor NOR3_42(g11773,g9400,g9479,g9603);
  nor NOR3_43(g11780,g9440,g9519,g9630);
  nor NOR3_44(g11781,g9442,g9522,g9633);
  nor NOR3_45(g11784,g9463,g9581,g9660);
  nor NOR3_46(g11785,g9464,g9583,g9663);
  nor NOR3_47(g11789,g9480,g9604,g9722);
  nor NOR3_48(g11790,g9497,g9621,g9745);
  nor NOR3_49(g11799,g9520,g9631,g9759);
  nor NOR3_50(g11800,g9523,g9634,g9762);
  nor NOR3_51(g11806,g9582,g9661,g9776);
  nor NOR3_52(g11807,g9584,g9664,g9779);
  nor NOR3_53(g11810,g9605,g9723,g9806);
  nor NOR3_54(g11811,g9606,g9725,g9809);
  nor NOR3_55(g11815,g9622,g9746,g9868);
  nor NOR3_56(g11822,g9632,g9760,g9888);
  nor NOR3_57(g11823,g9635,g9763,g9891);
  nor NOR3_58(g11828,g9639,g9764,g9892);
  nor NOR3_59(g11830,g9647,g9773,g9901);
  nor NOR3_60(g11831,g9648,g9775,g9904);
  nor NOR3_61(g11832,g9662,g9777,g9905);
  nor NOR3_62(g11833,g9665,g9780,g9908);
  nor NOR3_63(g11839,g9724,g9807,g9922);
  nor NOR3_64(g11840,g9726,g9810,g9925);
  nor NOR3_65(g11843,g9747,g9869,g9952);
  nor NOR3_66(g11844,g9748,g9871,g9955);
  nor NOR3_67(g11855,g9761,g9889,g10009);
  nor NOR3_68(g11860,g9765,g9893,g10012);
  nor NOR3_69(g11861,g9766,g9894,g10013);
  nor NOR3_70(g11863,g9774,g9902,g10035);
  nor NOR3_71(g11864,g9778,g9906,g10042);
  nor NOR3_72(g11865,g9781,g9909,g10045);
  nor NOR3_73(g11870,g9785,g9910,g10046);
  nor NOR3_74(g11872,g9793,g9919,g10055);
  nor NOR3_75(g11873,g9794,g9921,g10058);
  nor NOR3_76(g11874,g9808,g9923,g10059);
  nor NOR3_77(g11875,g9811,g9926,g10062);
  nor NOR3_78(g11881,g9870,g9953,g10076);
  nor NOR3_79(g11882,g9872,g9956,g10079);
  nor NOR3_80(g11889,g9887,g10007,g10101);
  nor NOR3_81(g11890,g9890,g10010,g10103);
  nor NOR3_82(g11896,g9903,g10036,g10112);
  nor NOR3_83(g11897,g9907,g10043,g10118);
  nor NOR3_84(g11902,g9911,g10047,g10121);
  nor NOR3_85(g11903,g9912,g10048,g10122);
  nor NOR3_86(g11905,g9920,g10056,g10144);
  nor NOR3_87(g11906,g9924,g10060,g10151);
  nor NOR3_88(g11907,g9927,g10063,g10154);
  nor NOR3_89(g11912,g9931,g10064,g10155);
  nor NOR3_90(g11914,g9939,g10073,g10164);
  nor NOR3_91(g11915,g9940,g10075,g10167);
  nor NOR3_92(g11916,g9954,g10077,g10168);
  nor NOR3_93(g11917,g9957,g10080,g10171);
  nor NOR3_94(g11928,g10008,g10102,g10192);
  nor NOR3_95(g11934,g10011,g10104,g10193);
  nor NOR3_96(g11935,g10014,g10106,g10196);
  nor NOR3_97(g11938,g10037,g10113,g10201);
  nor NOR3_98(g11939,g10041,g10116,g10206);
  nor NOR3_99(g11940,g10044,g10119,g10208);
  nor NOR3_100(g11946,g10057,g10145,g10217);
  nor NOR3_101(g11947,g10061,g10152,g10223);
  nor NOR3_102(g11952,g10065,g10156,g10226);
  nor NOR3_103(g11953,g10066,g10157,g10227);
  nor NOR3_104(g11955,g10074,g10165,g10249);
  nor NOR3_105(g11956,g10078,g10169,g10256);
  nor NOR3_106(g11957,g10081,g10172,g10259);
  nor NOR3_107(g11962,g10085,g10173,g10260);
  nor NOR3_108(g11964,g10093,g10182,g10269);
  nor NOR3_109(g11965,g10094,g10184,g10272);
  nor NOR3_110(g11974,g10105,g10194,g10279);
  nor NOR3_111(g11975,g10107,g10197,g10282);
  nor NOR3_112(g11979,g10114,g10202,g10288);
  nor NOR3_113(g11980,g10115,g10204,g10291);
  nor NOR3_114(g11981,g10117,g10207,g10294);
  nor NOR3_115(g11987,g10120,g10209,g10295);
  nor NOR3_116(g11988,g10123,g10211,g10298);
  nor NOR3_117(g11991,g10146,g10218,g10303);
  nor NOR3_118(g11992,g10150,g10221,g10308);
  nor NOR3_119(g11993,g10153,g10224,g10310);
  nor NOR3_120(g11999,g10166,g10250,g10319);
  nor NOR3_121(g12000,g10170,g10257,g10325);
  nor NOR3_122(g12005,g10174,g10261,g10328);
  nor NOR3_123(g12006,g10175,g10262,g10329);
  nor NOR3_124(g12008,g10183,g10270,g10351);
  nor NOR3_125(g12026,g10195,g10280,g10360);
  nor NOR3_126(g12033,g10199,g10284,g10362);
  nor NOR3_127(g12034,g10200,g10286,g10365);
  nor NOR3_128(g12035,g10203,g10289,g10367);
  nor NOR3_129(g12036,g10205,g10292,g10370);
  nor NOR3_130(g12043,g10210,g10296,g10372);
  nor NOR3_131(g12044,g10212,g10299,g10375);
  nor NOR3_132(g12048,g10219,g10304,g10381);
  nor NOR3_133(g12049,g10220,g10306,g10384);
  nor NOR3_134(g12050,g10222,g10309,g10387);
  nor NOR3_135(g12056,g10225,g10311,g10388);
  nor NOR3_136(g12057,g10228,g10313,g10391);
  nor NOR3_137(g12060,g10251,g10320,g10396);
  nor NOR3_138(g12061,g10255,g10323,g10401);
  nor NOR3_139(g12062,g10258,g10326,g10403);
  nor NOR3_140(g12068,g10271,g10352,g10412);
  nor NOR3_141(g12079,g10281,g10361,g10422);
  nor NOR3_142(g12080,g10285,g10363,g10430);
  nor NOR3_143(g12081,g10287,g10366,g10433);
  nor NOR3_144(g12082,g10290,g10368,g10435);
  nor NOR3_145(g12083,g10293,g10371,g10438);
  nor NOR3_146(g12090,g10297,g10373,g10439);
  nor NOR3_147(g12097,g10301,g10377,g10441);
  nor NOR3_148(g12098,g10302,g10379,g10444);
  nor NOR3_149(g12099,g10305,g10382,g10446);
  nor NOR3_150(g12100,g10307,g10385,g10449);
  nor NOR3_151(g12107,g10312,g10389,g10451);
  nor NOR3_152(g12108,g10314,g10392,g10454);
  nor NOR3_153(g12112,g10321,g10397,g10460);
  nor NOR3_154(g12113,g10322,g10399,g10463);
  nor NOR3_155(g12114,g10324,g10402,g10466);
  nor NOR3_156(g12120,g10327,g10404,g10467);
  nor NOR3_157(g12121,g10330,g10406,g10470);
  nor NOR3_158(g12124,g10353,g10413,g10475);
  nor NOR3_159(g12145,g10364,g10431,g10492);
  nor NOR3_160(g12146,g10369,g10436,g10496);
  nor NOR3_161(g12151,g10374,g10440,g10498);
  nor NOR3_162(g12152,g10378,g10442,g10506);
  nor NOR3_163(g12153,g10380,g10445,g10509);
  nor NOR3_164(g12154,g10383,g10447,g10511);
  nor NOR3_165(g12155,g10386,g10450,g10514);
  nor NOR3_166(g12162,g10390,g10452,g10515);
  nor NOR3_167(g12169,g10394,g10456,g10517);
  nor NOR3_168(g12170,g10395,g10458,g10520);
  nor NOR3_169(g12171,g10398,g10461,g10522);
  nor NOR3_170(g12172,g10400,g10464,g10525);
  nor NOR3_171(g12179,g10405,g10468,g10527);
  nor NOR3_172(g12180,g10407,g10471,g10530);
  nor NOR3_173(g12184,g10414,g10476,g10536);
  nor NOR3_174(g12185,g10415,g10478,g10539);
  nor NOR3_175(g12192,g10423,g10485,g10548);
  nor NOR3_176(g12193,g10432,g10493,g10555);
  nor NOR3_177(g12194,g10434,g10494,g10556);
  nor NOR3_178(g12195,g10437,g10497,g10558);
  nor NOR3_179(g12207,g10443,g10507,g10566);
  nor NOR3_180(g12208,g10448,g10512,g10570);
  nor NOR3_181(g12213,g10453,g10516,g10572);
  nor NOR3_182(g12214,g10457,g10518,g10580);
  nor NOR3_183(g12215,g10459,g10521,g10583);
  nor NOR3_184(g12216,g10462,g10523,g10585);
  nor NOR3_185(g12217,g10465,g10526,g10588);
  nor NOR3_186(g12224,g10469,g10528,g10589);
  nor NOR3_187(g12231,g10473,g10532,g10591);
  nor NOR3_188(g12232,g10474,g10534,g10594);
  nor NOR3_189(g12233,g10477,g10537,g10596);
  nor NOR3_190(g12234,g10479,g10540,g10599);
  nor NOR3_191(g12245,g10495,g10557,g10604);
  nor NOR3_192(g12247,g10499,g10559,g10605);
  nor NOR3_193(g12248,g10508,g10567,g10612);
  nor NOR3_194(g12249,g10510,g10568,g10613);
  nor NOR3_195(g12250,g10513,g10571,g10615);
  nor NOR3_196(g12262,g10519,g10581,g10623);
  nor NOR3_197(g12263,g10524,g10586,g10627);
  nor NOR3_198(g12268,g10529,g10590,g10629);
  nor NOR3_199(g12269,g10533,g10592,g10637);
  nor NOR3_200(g12270,g10535,g10595,g10640);
  nor NOR3_201(g12271,g10538,g10597,g10642);
  nor NOR3_202(g12272,g10541,g10600,g10645);
  nor NOR3_203(g12288,g10569,g10614,g10651);
  nor NOR3_204(g12290,g10573,g10616,g10652);
  nor NOR3_205(g12291,g10582,g10624,g10659);
  nor NOR3_206(g12292,g10584,g10625,g10660);
  nor NOR3_207(g12293,g10587,g10628,g10662);
  nor NOR3_208(g12305,g10593,g10638,g10670);
  nor NOR3_209(g12306,g10598,g10643,g10674);
  nor NOR3_210(g12324,g10626,g10661,g10681);
  nor NOR3_211(g12326,g10630,g10663,g10682);
  nor NOR3_212(g12327,g10639,g10671,g10689);
  nor NOR3_213(g12328,g10641,g10672,g10690);
  nor NOR3_214(g12329,g10644,g10675,g10692);
  nor NOR3_215(g12339,g10650,g10678,g10704);
  nor NOR3_216(g12352,g10673,g10691,g10710);
  nor NOR3_217(g12369,g10680,g10707,g10724);
  nor NOR3_218(g12388,g10709,g10727,g10745);
  nor NOR3_219(g12418,g10729,g10748,g10764);
  nor NOR2_2(g12431,g8580,g10730);
  nor NOR2_3(g12436,g8587,g10749);
  nor NOR2_4(g12441,g8594,g10767);
  nor NOR2_5(g12446,g8605,g10773);
  nor NOR2_6(g12451,g499,g8983);
  nor NOR3_220(g12457,g9009,g9033,g9048);
  nor NOR3_221(g12467,g9034,g9056,g9065);
  nor NOR3_222(g12482,g9057,g9073,g9082);
  nor NOR3_223(g12487,g10108,g10198,g10283);
  nor NOR3_224(g12499,g9074,g9090,g9101);
  nor NOR3_225(g12507,g10213,g10300,g10376);
  nor NOR3_226(g12524,g10315,g10393,g10455);
  nor NOR3_227(g12539,g10408,g10472,g10531);
  nor NOR3_228(g12698,g11347,g11420,g8327);
  nor NOR3_229(g12747,g11421,g8328,g8385);
  nor NOR3_230(g12755,g11431,g8339,g8394);
  nor NOR2_7(g12780,g9187,g9161);
  nor NOR3_231(g12781,g8329,g8386,g8431);
  nor NOR3_232(g12789,g8340,g8395,g8437);
  nor NOR3_233(g12797,g8350,g8406,g8446);
  nor NOR3_234(g12814,g8387,g8432,g8463);
  nor NOR2_8(g12819,g9248,g9203);
  nor NOR3_235(g12820,g8396,g8438,g8466);
  nor NOR3_236(g12828,g8407,g8447,g8472);
  nor NOR3_237(g12836,g8417,g8458,g8481);
  nor NOR3_238(g12849,g8433,g8464,g8485);
  nor NOR3_239(g12852,g8439,g8467,g8488);
  nor NOR2_9(g12857,g9326,g9264);
  nor NOR3_240(g12858,g8448,g8473,g8491);
  nor NOR3_241(g12866,g8459,g8482,g8497);
  nor NOR3_242(g12880,g8465,g8486,g8502);
  nor NOR2_10(g12883,g10038,g6284);
  nor NOR3_243(g12890,g8468,g8489,g8505);
  nor NOR3_244(g12893,g8474,g8492,g8508);
  nor NOR2_11(g12898,g9407,g9342);
  nor NOR3_245(g12899,g8483,g8498,g8511);
  nor NOR3_246(g12912,g8484,g8500,g8515);
  nor NOR3_247(g12913,g8487,g8503,g8518);
  nor NOR3_248(g12920,g8490,g8506,g8521);
  nor NOR2_12(g12923,g10147,g6421);
  nor NOR3_249(g12930,g8493,g8509,g8524);
  nor NOR3_250(g12933,g8499,g8512,g8527);
  nor NOR3_251(g12939,g8501,g8516,g8531);
  nor NOR3_252(g12941,g8504,g8519,g8534);
  nor NOR3_253(g12942,g8507,g8522,g8537);
  nor NOR3_254(g12949,g8510,g8525,g8540);
  nor NOR2_13(g12952,g10252,g6626);
  nor NOR3_255(g12959,g8513,g8528,g8543);
  nor NOR3_256(g12967,g8517,g8532,g8546);
  nor NOR3_257(g12968,g8520,g8535,g8548);
  nor NOR3_258(g12970,g8523,g8538,g8551);
  nor NOR3_259(g12971,g8526,g8541,g8554);
  nor NOR3_260(g12978,g8529,g8544,g8557);
  nor NOR2_14(g12981,g10354,g6890);
  nor NOR3_261(g12991,g8536,g8549,g8559);
  nor NOR3_262(g12992,g8539,g8552,g8561);
  nor NOR3_263(g12994,g8542,g8555,g8564);
  nor NOR3_264(g12995,g8545,g8558,g8567);
  nor NOR3_265(g13001,g8553,g8562,g8570);
  nor NOR3_266(g13002,g8556,g8565,g8572);
  nor NOR3_267(g13022,g8566,g8573,g8576);
  nor NOR4_4(g13024,g11481,g8045,g7928,g7880);
  nor NOR3_268(g13111,g8601,g8612,g8621);
  nor NOR3_269(g13124,g8613,g8625,g8631);
  nor NOR3_270(g13135,g8626,g8635,g8650);
  nor NOR3_271(g13143,g8636,g8654,g8666);
  nor NOR3_272(g13149,g8676,g8687,g8703);
  nor NOR3_273(g13155,g8688,g8705,g8722);
  nor NOR3_274(g13160,g8704,g8717,g8751);
  nor NOR3_275(g13164,g8706,g8724,g8760);
  nor NOR3_276(g13171,g8723,g8755,g8774);
  nor NOR3_277(g13175,g8725,g8762,g8783);
  nor NOR3_278(g13182,g8761,g8778,g8797);
  nor NOR3_279(g13194,g8784,g8801,g8816);
  nor NOR3_280(g13228,g8841,g8861,g8892);
  nor NOR3_281(g13251,g8868,g8899,g8932);
  nor NOR3_282(g13274,g8906,g8939,g8972);
  nor NOR4_5(g13286,g11481,g11332,g11190,g7880);
  nor NOR3_283(g13299,g8946,g8979,g9004);
  nor NOR4_6(g13310,g11481,g11332,g11190,g11069);
  nor NOR4_7(g13313,g8183,g11332,g11190,g7880);
  nor NOR4_8(g13331,g8183,g11332,g11190,g11069);
  nor NOR4_9(g13332,g11481,g8045,g11190,g7880);
  nor NOR4_10(g13353,g11481,g8045,g11190,g11069);
  nor NOR4_11(g13354,g8183,g8045,g11190,g7880);
  nor NOR4_12(g13374,g8183,g8045,g11190,g11069);
  nor NOR4_13(g13375,g11481,g11332,g7928,g7880);
  nor NOR3_284(g13378,g9026,g9047,g9061);
  nor NOR4_14(g13401,g11481,g11332,g7928,g11069);
  nor NOR4_15(g13404,g8183,g11332,g7928,g7880);
  nor NOR2_15(g15661,g11737,g7345);
  nor NOR2_16(g15797,g13305,g7143);
  nor NOR2_17(g15873,g11617,g7562);
  nor NOR2_18(g15959,g2814,g13082);
  nor NOR2_19(g15978,g11737,g7152);
  nor NOR3_285(g16020,g6200,g12457,g10952);
  nor NOR3_286(g16036,g6289,g12467,g10952);
  nor NOR3_287(g16058,g6426,g12482,g10952);
  nor NOR3_288(g16082,g10952,g6140,g12487);
  nor NOR3_289(g16094,g6631,g12499,g10952);
  nor NOR3_290(g16120,g10952,g6161,g12507);
  nor NOR3_291(g16171,g10952,g6188,g12524);
  nor NOR3_292(g16230,g10952,g6220,g12539);
  nor NOR2_20(g16498,g14158,g14347);
  nor NOR2_21(g16520,g14273,g14459);
  nor NOR2_22(g16551,g14395,g14546);
  nor NOR3_293(g16567,g15904,g15880,g15859);
  nor NOR3_294(g16570,g15904,g15880,g14630);
  nor NOR2_23(g16583,g14507,g14601);
  nor NOR3_295(g16591,g15933,g15913,g15890);
  nor NOR3_296(g16594,g15933,g15913,g14650);
  nor NOR3_297(g16611,g15962,g15942,g15923);
  nor NOR3_298(g16614,g15962,g15942,g14677);
  nor NOR3_299(g16629,g15981,g15971,g15952);
  nor NOR3_300(g16632,g15981,g15971,g14711);
  nor NOR3_301(g16643,g15904,g14642,g15859);
  nor NOR2_24(g16654,g14690,g12477);
  nor NOR3_302(g16655,g15933,g14669,g15890);
  nor NOR2_25(g16671,g14724,g12494);
  nor NOR3_303(g16672,g15962,g14703,g15923);
  nor NOR2_26(g16679,g14797,g14895);
  nor NOR2_27(g16692,g14752,g12514);
  nor NOR3_304(g16693,g15981,g14737,g15952);
  nor NOR2_28(g16705,g14849,g14976);
  nor NOR2_29(g16718,g14773,g12531);
  nor NOR2_30(g16736,g14922,g15065);
  nor NOR2_31(g16778,g15003,g15161);
  nor NOR2_32(g16802,g13469,g3897);
  nor NOR2_33(g16803,g15593,g12908);
  nor NOR2_34(g16823,g5362,g13469);
  nor NOR2_35(g16824,g15658,g12938);
  nor NOR2_36(g16829,g14956,g12564);
  nor NOR2_37(g16835,g15717,g12966);
  nor NOR2_38(g16841,g15021,g12607);
  nor NOR2_39(g16844,g15754,g12989);
  nor NOR2_40(g16845,g15755,g12990);
  nor NOR2_41(g16847,g15095,g12650);
  nor NOR2_42(g16851,g15781,g13000);
  nor NOR2_43(g16853,g15801,g13009);
  nor NOR2_44(g16854,g15802,g13010);
  nor NOR2_45(g16857,g15817,g13023);
  nor NOR2_46(g16860,g15828,g13031);
  nor NOR2_47(g16861,g15829,g13032);
  nor NOR2_48(g16866,g15840,g13042);
  nor NOR2_49(g16880,g15852,g13056);
  nor NOR3_305(g17012,g14657,g14642,g15859);
  nor NOR3_306(g17025,g15904,g15880,g15859);
  nor NOR3_307(g17042,g14691,g14669,g15890);
  nor NOR3_308(g17051,g14657,g15880,g14630);
  nor NOR3_309(g17059,g15933,g15913,g15890);
  nor NOR3_310(g17076,g14725,g14703,g15923);
  nor NOR3_311(g17086,g14691,g15913,g14650);
  nor NOR3_312(g17094,g15962,g15942,g15923);
  nor NOR3_313(g17111,g14753,g14737,g15952);
  nor NOR3_314(g17124,g14725,g15942,g14677);
  nor NOR3_315(g17132,g15981,g15971,g15952);
  nor NOR3_316(g17151,g14753,g15971,g14711);
  nor NOR2_50(g17186,g7949,g14144);
  nor NOR2_51(g17197,g8000,g14259);
  nor NOR2_52(g17204,g8075,g14381);
  nor NOR2_53(g17209,g8160,g14493);
  nor NOR2_54(g17213,g4326,g14442);
  nor NOR2_55(g17215,g15904,g14642);
  nor NOR2_56(g17216,g4495,g14529);
  nor NOR2_57(g17218,g15933,g14669);
  nor NOR2_58(g17219,g4671,g14584);
  nor NOR2_59(g17220,g15962,g14703);
  nor NOR2_60(g17221,g4848,g14618);
  nor NOR2_61(g17222,g15998,g16003);
  nor NOR2_62(g17223,g15981,g14737);
  nor NOR2_63(g17224,g16004,g16009);
  nor NOR2_64(g17225,g16008,g16015);
  nor NOR2_65(g17226,g16010,g16017);
  nor NOR2_66(g17228,g16016,g16029);
  nor NOR2_67(g17229,g16019,g16032);
  nor NOR2_68(g17234,g16028,g16045);
  nor NOR2_69(g17235,g16030,g16047);
  nor NOR2_70(g17236,g16033,g16051);
  nor NOR2_71(g17246,g16046,g16066);
  nor NOR2_72(g17247,g16050,g16070);
  nor NOR2_73(g17248,g16052,g16072);
  nor NOR2_74(g17269,g16067,g16100);
  nor NOR2_75(g17270,g16071,g16104);
  nor NOR2_76(g17271,g16073,g16106);
  nor NOR2_77(g17302,g16103,g16135);
  nor NOR2_78(g17303,g16105,g16137);
  nor NOR2_79(g17340,g16136,g16183);
  nor NOR2_80(g17341,g16138,g16185);
  nor NOR2_81(g17383,g16184,g16238);
  nor NOR2_82(g17429,g16239,g16288);
  nor NOR2_83(g17507,g16298,g13318);
  nor NOR2_84(g17896,g14352,g16020);
  nor NOR2_85(g18007,g14464,g16036);
  nor NOR2_86(g18085,g16085,g6363);
  nor NOR2_87(g18124,g14551,g16058);
  nor NOR2_88(g18201,g16123,g6568);
  nor NOR2_89(g18240,g14606,g16094);
  nor NOR2_90(g18308,g16174,g6832);
  nor NOR2_91(g18352,g16082,g14249);
  nor NOR2_92(g18401,g16233,g7134);
  nor NOR2_93(g18430,g16020,g14352);
  nor NOR2_94(g18447,g16120,g14371);
  nor NOR2_95(g18503,g16036,g14464);
  nor NOR2_96(g18520,g16171,g14483);
  nor NOR2_97(g18548,g14249,g16082);
  nor NOR2_98(g18567,g16058,g14551);
  nor NOR2_99(g18584,g16230,g14570);
  nor NOR2_100(g18590,g16439,g7522);
  nor NOR2_101(g18598,g14371,g16120);
  nor NOR2_102(g18617,g16094,g14606);
  nor NOR2_103(g18623,g15902,g2814);
  nor NOR2_104(g18626,g16463,g7549);
  nor NOR2_105(g18630,g14483,g16171);
  nor NOR2_106(g18639,g14570,g16230);
  nor NOR2_107(g18669,g13623,g13634);
  nor NOR2_108(g18678,g13625,g11771);
  nor NOR2_109(g18707,g13636,g11788);
  nor NOR2_110(g18719,g13643,g13656);
  nor NOR2_111(g18726,g13645,g11805);
  nor NOR2_112(g18743,g13648,g11814);
  nor NOR2_113(g18754,g13655,g11816);
  nor NOR2_114(g18755,g13871,g12274);
  nor NOR2_115(g18763,g13671,g11838);
  nor NOR2_116(g18780,g13674,g11847);
  nor NOR2_117(g18781,g13675,g11851);
  nor NOR2_118(g18782,g13676,g13705);
  nor NOR2_119(g18794,g13701,g11880);
  nor NOR2_120(g18803,g13704,g11885);
  nor NOR2_121(g18804,g13905,g12331);
  nor NOR2_122(g18820,g13738,g11922);
  nor NOR2_123(g18821,g13740,g11926);
  nor NOR2_124(g18835,g13788,g11966);
  nor NOR2_125(g18836,g13789,g11967);
  nor NOR2_126(g18837,g13998,g12376);
  nor NOR2_127(g18852,g13815,g12012);
  nor NOR2_128(g18866,g13834,g12069);
  nor NOR2_129(g18867,g13835,g12070);
  nor NOR2_130(g18868,g14143,g12419);
  nor NOR2_131(g18883,g13846,g12128);
  nor NOR2_132(g18885,g13847,g12129);
  nor NOR2_133(g18906,g13855,g12186);
  nor NOR2_134(g18907,g14336,g12429);
  nor NOR2_135(g18942,g13870,g12273);
  nor NOR2_136(g18957,g13884,g12307);
  nor NOR2_137(g18968,g13904,g12330);
  nor NOR2_138(g18975,g13944,g12353);
  nor NOR2_139(g19144,g17268,g14884);
  nor NOR2_140(g19149,g17339,g15020);
  nor NOR2_141(g19153,g17381,g15093);
  nor NOR2_142(g19154,g17382,g15094);
  nor NOR2_143(g19157,g17428,g15171);
  nor NOR2_144(g19160,g17446,g15178);
  nor NOR2_145(g19162,g17485,g15243);
  nor NOR2_146(g19163,g17486,g15244);
  nor NOR2_147(g19165,g17526,g15264);
  nor NOR2_148(g19167,g17556,g15320);
  nor NOR2_149(g19171,g17616,g15356);
  nor NOR2_150(g19172,g17635,g15388);
  nor NOR2_151(g19173,g17636,g15389);
  nor NOR2_152(g19177,g17713,g15442);
  nor NOR2_153(g19178,g17718,g15452);
  nor NOR2_154(g19179,g17719,g15453);
  nor NOR2_155(g19184,g17798,g15520);
  nor NOR2_156(g19219,g18165,g15753);
  nor NOR2_157(g20008,g18977,g7338);
  nor NOR2_158(g20054,g19001,g16867);
  nor NOR2_159(g20095,g16507,g16895);
  nor NOR2_160(g20120,g16529,g16924);
  nor NOR2_161(g20150,g16560,g16954);
  nor NOR2_162(g20153,g16536,g7583);
  nor NOR2_163(g20299,g16665,g16884);
  nor NOR2_164(g20310,g16850,g13654);
  nor NOR2_165(g20314,g13646,g16855);
  nor NOR2_166(g20318,g16686,g16913);
  nor NOR2_167(g20333,g13672,g16859);
  nor NOR2_168(g20337,g16712,g16943);
  nor NOR2_169(g20343,g16856,g13703);
  nor NOR2_170(g20353,g13702,g16864);
  nor NOR2_171(g20357,g16743,g16974);
  nor NOR2_172(g20375,g13739,g16879);
  nor NOR2_173(g20376,g16865,g13787);
  nor NOR2_174(g20417,g16907,g13833);
  nor NOR2_175(g20682,g19160,g10024);
  nor NOR2_176(g20717,g19165,g10133);
  nor NOR2_177(g20752,g19171,g10238);
  nor NOR2_178(g20789,g19177,g10340);
  nor NOR2_179(g20841,g14767,g19552);
  nor NOR2_180(g20874,g17301,g19594);
  nor NOR2_181(g20875,g19584,g17352);
  nor NOR2_182(g20876,g19585,g17353);
  nor NOR2_183(g20877,g3919,g19830);
  nor NOR2_184(g20878,g19600,g17395);
  nor NOR2_185(g20879,g19601,g17396);
  nor NOR2_186(g20880,g19602,g17397);
  nor NOR2_187(g20881,g19603,g17398);
  nor NOR2_188(g20882,g19614,g17408);
  nor NOR2_189(g20883,g19615,g17409);
  nor NOR2_190(g20884,g5394,g19830);
  nor NOR2_191(g20891,g19626,g17447);
  nor NOR2_192(g20892,g19627,g17448);
  nor NOR2_193(g20893,g19628,g17449);
  nor NOR2_194(g20894,g19629,g17450);
  nor NOR2_195(g20895,g19633,g17461);
  nor NOR2_196(g20896,g19634,g17462);
  nor NOR2_197(g20897,g19635,g17463);
  nor NOR2_198(g20898,g19636,g17464);
  nor NOR2_199(g20899,g19647,g17474);
  nor NOR2_200(g20900,g19648,g17475);
  nor NOR2_201(g20901,g19660,g17508);
  nor NOR2_202(g20902,g19661,g17509);
  nor NOR2_203(g20903,g19662,g17510);
  nor NOR2_204(g20910,g19666,g17527);
  nor NOR2_205(g20911,g19667,g17528);
  nor NOR2_206(g20912,g19668,g17529);
  nor NOR2_207(g20913,g19669,g17530);
  nor NOR2_208(g20914,g19673,g17541);
  nor NOR2_209(g20915,g19674,g17542);
  nor NOR2_210(g20916,g19675,g17543);
  nor NOR2_211(g20917,g19676,g17544);
  nor NOR2_212(g20918,g19687,g17554);
  nor NOR2_213(g20919,g19688,g17555);
  nor NOR2_214(g20920,g19691,g19726);
  nor NOR2_215(g20921,g19697,g17576);
  nor NOR2_216(g20922,g19698,g17577);
  nor NOR2_217(g20923,g19699,g17578);
  nor NOR2_218(g20924,g19700,g15257);
  nor NOR2_219(g20925,g19708,g17598);
  nor NOR2_220(g20926,g19709,g17599);
  nor NOR2_221(g20927,g19710,g17600);
  nor NOR2_222(g20934,g19714,g17617);
  nor NOR2_223(g20935,g19715,g17618);
  nor NOR2_224(g20936,g19716,g17619);
  nor NOR2_225(g20937,g19717,g17620);
  nor NOR2_226(g20938,g19721,g17631);
  nor NOR2_227(g20939,g19722,g17632);
  nor NOR2_228(g20940,g19723,g17633);
  nor NOR2_229(g20941,g19724,g17634);
  nor NOR2_230(g20944,g19731,g17652);
  nor NOR2_231(g20945,g19732,g17653);
  nor NOR2_232(g20946,g19733,g17654);
  nor NOR2_233(g20947,g19734,g15335);
  nor NOR2_234(g20948,g19735,g15336);
  nor NOR2_235(g20949,g19741,g17673);
  nor NOR2_236(g20950,g19742,g17674);
  nor NOR2_237(g20951,g19743,g17675);
  nor NOR2_238(g20952,g19744,g15349);
  nor NOR2_239(g20953,g19752,g17695);
  nor NOR2_240(g20954,g19753,g17696);
  nor NOR2_241(g20955,g19754,g17697);
  nor NOR2_242(g20962,g19758,g17714);
  nor NOR2_243(g20963,g19759,g17715);
  nor NOR2_244(g20964,g19760,g17716);
  nor NOR2_245(g20965,g19761,g17717);
  nor NOR2_246(g20966,g19765,g17734);
  nor NOR2_247(g20967,g19766,g17735);
  nor NOR2_248(g20968,g19767,g17736);
  nor NOR2_249(g20969,g19768,g15402);
  nor NOR2_250(g20970,g19769,g15403);
  nor NOR2_251(g20972,g19774,g17752);
  nor NOR2_252(g20973,g19775,g17753);
  nor NOR2_253(g20974,g19776,g17754);
  nor NOR2_254(g20975,g19777,g15421);
  nor NOR2_255(g20976,g19778,g15422);
  nor NOR2_256(g20977,g19784,g17773);
  nor NOR2_257(g20978,g19785,g17774);
  nor NOR2_258(g20979,g19786,g17775);
  nor NOR2_259(g20980,g19787,g15435);
  nor NOR2_260(g20981,g19795,g17795);
  nor NOR2_261(g20982,g19796,g17796);
  nor NOR2_262(g20983,g19797,g17797);
  nor NOR2_263(g20989,g19802,g17812);
  nor NOR2_264(g20990,g19803,g17813);
  nor NOR2_265(g20991,g19804,g17814);
  nor NOR2_266(g20992,g19805,g15470);
  nor NOR2_267(g20993,g19807,g17835);
  nor NOR2_268(g20994,g19808,g17836);
  nor NOR2_269(g20995,g19809,g17837);
  nor NOR2_270(g20996,g19810,g15486);
  nor NOR2_271(g20997,g19811,g15487);
  nor NOR2_272(g20999,g19816,g17853);
  nor NOR2_273(g21000,g19817,g17854);
  nor NOR2_274(g21001,g19818,g17855);
  nor NOR2_275(g21002,g19819,g15505);
  nor NOR2_276(g21003,g19820,g15506);
  nor NOR2_277(g21004,g19826,g17874);
  nor NOR2_278(g21005,g19827,g17875);
  nor NOR2_279(g21006,g19828,g17876);
  nor NOR2_280(g21007,g19829,g15519);
  nor NOR2_281(g21008,g19836,g17877);
  nor NOR2_282(g21009,g19839,g17900);
  nor NOR2_283(g21010,g19840,g17901);
  nor NOR2_284(g21011,g19841,g17902);
  nor NOR2_285(g21015,g19846,g17924);
  nor NOR2_286(g21016,g19847,g17925);
  nor NOR2_287(g21017,g19848,g17926);
  nor NOR2_288(g21018,g19849,g15556);
  nor NOR2_289(g21019,g19851,g17947);
  nor NOR2_290(g21020,g19852,g17948);
  nor NOR2_291(g21021,g19853,g17949);
  nor NOR2_292(g21022,g19854,g15572);
  nor NOR2_293(g21023,g19855,g15573);
  nor NOR2_294(g21025,g19860,g17965);
  nor NOR2_295(g21026,g19861,g17966);
  nor NOR2_296(g21027,g19862,g17967);
  nor NOR2_297(g21028,g19863,g15591);
  nor NOR2_298(g21029,g19864,g15592);
  nor NOR2_299(g21031,g19869,g17989);
  nor NOR2_300(g21032,g19870,g17990);
  nor NOR2_301(g21033,g19872,g18011);
  nor NOR2_302(g21034,g19873,g18012);
  nor NOR2_303(g21035,g19874,g18013);
  nor NOR2_304(g21039,g19879,g18035);
  nor NOR2_305(g21040,g19880,g18036);
  nor NOR2_306(g21041,g19881,g18037);
  nor NOR2_307(g21042,g19882,g15634);
  nor NOR2_308(g21043,g19884,g18058);
  nor NOR2_309(g21044,g19885,g18059);
  nor NOR2_310(g21045,g19886,g18060);
  nor NOR2_311(g21046,g19887,g15650);
  nor NOR2_312(g21047,g19888,g15651);
  nor NOR2_313(g21048,g19889,g18062);
  nor NOR2_314(g21051,g19895,g18088);
  nor NOR2_315(g21052,g19900,g18106);
  nor NOR2_316(g21053,g19901,g18107);
  nor NOR2_317(g21054,g19903,g18128);
  nor NOR2_318(g21055,g19904,g18129);
  nor NOR2_319(g21056,g19905,g18130);
  nor NOR2_320(g21060,g19910,g18152);
  nor NOR2_321(g21061,g19911,g18153);
  nor NOR2_322(g21062,g19912,g18154);
  nor NOR2_323(g21063,g19913,g15710);
  nor NOR2_324(g21065,g19914,g18169);
  nor NOR2_325(g21070,g19920,g18204);
  nor NOR2_326(g21071,g19925,g18222);
  nor NOR2_327(g21072,g19926,g18223);
  nor NOR2_328(g21073,g19928,g18244);
  nor NOR2_329(g21074,g19929,g18245);
  nor NOR2_330(g21075,g19930,g18246);
  nor NOR2_331(g21080,g19935,g18311);
  nor NOR2_332(g21081,g19940,g18329);
  nor NOR2_333(g21082,g19941,g18330);
  nor NOR2_334(g21083,g19943,g18333);
  nor NOR2_335(g21084,g20011,g20048);
  nor NOR2_336(g21094,g19952,g18404);
  nor NOR3_317(g21095,g20012,g20049,g20084);
  nor NOR3_318(g21096,g20013,g20051,g20087);
  nor NOR3_319(g21104,g20050,g20085,g20106);
  nor NOR3_320(g21105,g20052,g20088,g20109);
  nor NOR3_321(g21106,g20053,g20090,g20112);
  nor NOR3_322(g21116,g20086,g20107,g20131);
  nor NOR3_323(g21117,g20089,g20110,g20133);
  nor NOR3_324(g21118,g20091,g20113,g20136);
  nor NOR3_325(g21119,g20092,g20115,g20139);
  nor NOR3_326(g21133,g20108,g20132,g20156);
  nor NOR3_327(g21134,g20111,g20134,g20157);
  nor NOR3_328(g21135,g20114,g20137,g20160);
  nor NOR3_329(g21147,g20135,g20158,g20188);
  nor NOR3_330(g21148,g20138,g20161,g20190);
  nor NOR2_337(g21149,g20015,g19981);
  nor NOR2_338(g21167,g20159,g20189);
  nor NOR3_331(g21168,g20162,g20191,g20220);
  nor NOR2_339(g21169,g20057,g20019);
  nor NOR2_340(g21183,g20192,g20221);
  nor NOR2_341(g21189,g20098,g20061);
  nor NOR2_342(g21204,g20123,g20102);
  nor NOR2_343(g21211,g19240,g19230);
  nor NOR2_344(g21219,g19253,g19243);
  nor NOR3_332(g21227,g18414,g18485,g20295);
  nor NOR2_345(g21228,g19388,g17118);
  nor NOR2_346(g21230,g19266,g19256);
  nor NOR2_347(g21233,g19418,g17145);
  nor NOR2_348(g21235,g19281,g19269);
  nor NOR2_349(g21238,g19954,g5890);
  nor NOR2_350(g21242,g19455,g17168);
  nor NOR2_351(g21246,g19984,g5929);
  nor NOR2_352(g21250,g19482,g17183);
  nor NOR2_353(g21255,g20022,g5963);
  nor NOR2_354(g21263,g20064,g5992);
  nor NOR2_355(g21316,g20460,g16111);
  nor NOR2_356(g21331,g20472,g16153);
  nor NOR2_357(g21346,g20480,g13247);
  nor NOR2_358(g21364,g20486,g13266);
  nor NOR2_359(g21385,g20492,g13289);
  nor NOR2_360(g21407,g20499,g13316);
  nor NOR2_361(g21432,g20502,g13335);
  nor NOR2_362(g21435,g20503,g16385);
  nor NOR2_363(g21467,g20506,g13355);
  nor NOR2_364(g21470,g20512,g16417);
  nor NOR2_365(g21502,g20525,g16445);
  nor NOR2_366(g21615,g16567,g19957);
  nor NOR3_333(g21618,g20016,g14079,g14165);
  nor NOR2_367(g21636,g20473,g6513);
  nor NOR2_368(g21643,g16591,g19987);
  nor NOR3_334(g21646,g20058,g14194,g14280);
  nor NOR2_369(g21665,g20507,g18352);
  nor NOR2_370(g21667,g20481,g6777);
  nor NOR2_371(g21674,g16611,g20025);
  nor NOR3_335(g21677,g20099,g14309,g14402);
  nor NOR2_372(g21694,g20526,g18447);
  nor NOR2_373(g21696,g20487,g7079);
  nor NOR2_374(g21703,g16629,g20067);
  nor NOR3_336(g21706,g20124,g14431,g14514);
  nor NOR2_375(g21711,g19830,g15780);
  nor NOR2_376(g21730,g20545,g18520);
  nor NOR2_377(g21732,g20493,g7329);
  nor NOR3_337(g21738,g19444,g17893,g14079);
  nor NOR2_378(g21739,g20507,g18430);
  nor NOR2_379(g21756,g19070,g18584);
  nor NOR3_338(g21762,g19471,g18004,g14194);
  nor NOR2_380(g21763,g20526,g18503);
  nor NOR3_339(g21778,g19494,g18121,g14309);
  nor NOR2_381(g21779,g20545,g18567);
  nor NOR3_340(g21793,g19515,g18237,g14431);
  nor NOR2_382(g21794,g19070,g18617);
  nor NOR2_383(g21796,g19830,g13004);
  nor NOR2_384(g21842,g13609,g19150);
  nor NOR2_385(g21843,g13619,g19155);
  nor NOR2_386(g21845,g13631,g19161);
  nor NOR2_387(g21847,g13642,g19166);
  nor NOR2_388(g21851,g19252,g8842);
  nor NOR2_389(g21878,g16964,g19228);
  nor NOR2_390(g21880,g13854,g19236);
  nor NOR2_391(g21882,g13862,g19248);
  nor NOR2_392(g21884,g19260,g19284);
  nor NOR2_393(g21887,g13519,g19289);
  nor NOR2_394(g21889,g19285,g19316);
  nor NOR2_395(g21890,g13530,g19307);
  nor NOR2_396(g21893,g13541,g19328);
  nor NOR2_397(g21894,g19317,g19356);
  nor NOR2_398(g21901,g13552,g19355);
  nor NOR2_399(g21968,g21234,g19476);
  nor NOR2_400(g21969,g20895,g10133);
  nor NOR2_401(g21970,g17182,g21226);
  nor NOR2_402(g21971,g21243,g19499);
  nor NOR2_403(g21972,g20914,g10238);
  nor NOR2_404(g21973,g21251,g19520);
  nor NOR2_405(g21974,g20938,g10340);
  nor NOR2_406(g21975,g21245,g21259);
  nor NOR3_341(g21980,g21252,g19531,g19540);
  nor NOR2_407(g21981,g21254,g21267);
  nor NOR3_342(g21987,g21260,g19541,g19544);
  nor NOR2_408(g21988,g21262,g21276);
  nor NOR3_343(g22000,g21268,g19545,g19547);
  nor NOR2_409(g22001,g21270,g21283);
  nor NOR3_344(g22013,g21277,g19548,g19551);
  nor NOR2_410(g22025,g21284,g19549);
  nor NOR2_411(g22026,g21083,g18407);
  nor NOR2_412(g22027,g21290,g19553);
  nor NOR2_413(g22028,g21291,g19554);
  nor NOR2_414(g22029,g21292,g19555);
  nor NOR2_415(g22030,g21298,g19557);
  nor NOR2_416(g22031,g21299,g19558);
  nor NOR2_417(g22032,g21300,g19559);
  nor NOR2_418(g22033,g21301,g19560);
  nor NOR2_419(g22034,g21302,g19561);
  nor NOR2_420(g22035,g21303,g19562);
  nor NOR2_421(g22037,g21304,g19564);
  nor NOR2_422(g22038,g21305,g19565);
  nor NOR2_423(g22039,g21306,g19566);
  nor NOR2_424(g22040,g21307,g19567);
  nor NOR2_425(g22041,g21308,g19568);
  nor NOR2_426(g22042,g21309,g19569);
  nor NOR2_427(g22043,g21310,g19570);
  nor NOR2_428(g22044,g21311,g19571);
  nor NOR2_429(g22045,g21312,g19572);
  nor NOR2_430(g22047,g21313,g19574);
  nor NOR2_431(g22048,g21314,g19575);
  nor NOR2_432(g22049,g21315,g19576);
  nor NOR2_433(g22054,g21319,g19586);
  nor NOR2_434(g22055,g21320,g19587);
  nor NOR2_435(g22056,g21321,g19588);
  nor NOR2_436(g22057,g21322,g19589);
  nor NOR2_437(g22058,g21323,g19590);
  nor NOR2_438(g22059,g21324,g19591);
  nor NOR2_439(g22060,g21325,g19592);
  nor NOR2_440(g22061,g21326,g19593);
  nor NOR2_441(g22063,g21328,g19597);
  nor NOR2_442(g22064,g21329,g19598);
  nor NOR2_443(g22065,g21330,g19599);
  nor NOR2_444(g22066,g21334,g19604);
  nor NOR2_445(g22067,g21335,g19605);
  nor NOR2_446(g22068,g21336,g19606);
  nor NOR2_447(g22073,g21337,g19616);
  nor NOR2_448(g22074,g21338,g19617);
  nor NOR2_449(g22075,g21339,g19618);
  nor NOR2_450(g22076,g21340,g19619);
  nor NOR2_451(g22077,g21341,g19620);
  nor NOR2_452(g22078,g21342,g19621);
  nor NOR2_453(g22079,g21343,g19623);
  nor NOR2_454(g22080,g21344,g19624);
  nor NOR2_455(g22081,g21345,g19625);
  nor NOR2_456(g22087,g21349,g19630);
  nor NOR2_457(g22088,g21350,g19631);
  nor NOR2_458(g22089,g21351,g19632);
  nor NOR2_459(g22090,g21352,g19637);
  nor NOR2_460(g22091,g21353,g19638);
  nor NOR2_461(g22092,g21354,g19639);
  nor NOR2_462(g22097,g21355,g19649);
  nor NOR2_463(g22098,g21356,g19650);
  nor NOR2_464(g22099,g21357,g19651);
  nor NOR2_465(g22100,g21360,g19653);
  nor NOR2_466(g22101,g21361,g19654);
  nor NOR2_467(g22102,g21362,g19655);
  nor NOR2_468(g22103,g21363,g19656);
  nor NOR2_469(g22104,g21367,g19663);
  nor NOR2_470(g22105,g21368,g19664);
  nor NOR2_471(g22106,g21369,g19665);
  nor NOR2_472(g22112,g21370,g19670);
  nor NOR2_473(g22113,g21371,g19671);
  nor NOR2_474(g22114,g21372,g19672);
  nor NOR2_475(g22115,g21373,g19677);
  nor NOR2_476(g22116,g21374,g19678);
  nor NOR2_477(g22117,g21375,g19679);
  nor NOR2_478(g22122,g21378,g19692);
  nor NOR2_479(g22123,g21379,g19693);
  nor NOR2_480(g22124,g21380,g19694);
  nor NOR2_481(g22125,g21381,g19695);
  nor NOR2_482(g22126,g21389,g19701);
  nor NOR2_483(g22127,g21390,g19702);
  nor NOR2_484(g22128,g21391,g19703);
  nor NOR2_485(g22129,g21392,g19704);
  nor NOR2_486(g22130,g21393,g19711);
  nor NOR2_487(g22131,g21394,g19712);
  nor NOR2_488(g22132,g21395,g19713);
  nor NOR2_489(g22138,g21396,g19718);
  nor NOR2_490(g22139,g21397,g19719);
  nor NOR2_491(g22140,g21398,g19720);
  nor NOR2_492(g22141,g21401,g19727);
  nor NOR2_493(g22142,g21402,g19728);
  nor NOR2_494(g22143,g21403,g19729);
  nor NOR2_495(g22144,g21410,g19730);
  nor NOR2_496(g22145,g21411,g19736);
  nor NOR2_497(g22146,g21412,g19737);
  nor NOR2_498(g22147,g21413,g19738);
  nor NOR2_499(g22148,g21414,g19739);
  nor NOR2_500(g22149,g21419,g19745);
  nor NOR2_501(g22150,g21420,g19746);
  nor NOR2_502(g22151,g21421,g19747);
  nor NOR2_503(g22152,g21422,g19748);
  nor NOR2_504(g22153,g21423,g19755);
  nor NOR2_505(g22154,g21424,g19756);
  nor NOR2_506(g22155,g21425,g19757);
  nor NOR2_507(g22161,g21428,g19764);
  nor NOR2_508(g22162,g21438,g19770);
  nor NOR2_509(g22163,g21439,g19771);
  nor NOR2_510(g22164,g21440,g19772);
  nor NOR2_511(g22165,g21444,g19773);
  nor NOR2_512(g22166,g21445,g19779);
  nor NOR2_513(g22167,g21446,g19780);
  nor NOR2_514(g22168,g21447,g19781);
  nor NOR2_515(g22169,g21448,g19782);
  nor NOR2_516(g22170,g21453,g19788);
  nor NOR2_517(g22171,g21454,g19789);
  nor NOR2_518(g22172,g21455,g19790);
  nor NOR2_519(g22173,g21456,g19791);
  nor NOR2_520(g22174,g19868,g21593);
  nor NOR2_521(g22177,g21476,g19806);
  nor NOR2_522(g22178,g21480,g19812);
  nor NOR2_523(g22179,g21481,g19813);
  nor NOR2_524(g22180,g21482,g19814);
  nor NOR2_525(g22181,g21486,g19815);
  nor NOR2_526(g22182,g21487,g19821);
  nor NOR2_527(g22183,g21488,g19822);
  nor NOR2_528(g22184,g21489,g19823);
  nor NOR2_529(g22185,g21490,g19824);
  nor NOR2_530(g22186,g21497,g19837);
  nor NOR2_531(g22189,g19899,g21622);
  nor NOR2_532(g22191,g21517,g19850);
  nor NOR2_533(g22192,g21521,g19856);
  nor NOR2_534(g22193,g21522,g19857);
  nor NOR2_535(g22194,g21523,g19858);
  nor NOR2_536(g22195,g21527,g19859);
  nor NOR2_537(g22198,g19924,g21650);
  nor NOR2_538(g22200,g21553,g19883);
  nor NOR2_539(g22204,g19939,g21681);
  nor NOR2_540(g22210,g21610,g19932);
  nor NOR2_541(g22216,g21635,g19944);
  nor NOR2_542(g22218,g21639,g19949);
  nor NOR2_543(g22227,g21658,g19953);
  nor NOR2_544(g22231,g21666,g19971);
  nor NOR2_545(g22234,g21670,g19976);
  nor NOR2_546(g22242,g21687,g19983);
  nor NOR2_547(g22247,g21695,g20001);
  nor NOR2_548(g22249,g21699,g20006);
  nor NOR2_549(g22263,g21723,g20021);
  nor NOR2_550(g22267,g21731,g20039);
  nor NOR2_551(g22269,g21735,g20044);
  nor NOR2_552(g22280,g21749,g20063);
  nor NOR2_553(g22284,g21757,g20081);
  nor NOR2_554(g22288,g20144,g21805);
  nor NOR2_555(g22299,g21773,g20104);
  nor NOR2_556(g22308,g20182,g21812);
  nor NOR2_557(g22336,g20216,g21818);
  nor NOR2_558(g22361,g20246,g21822);
  nor NOR2_559(g22454,g17012,g21891);
  nor NOR2_560(g22493,g17042,g21899);
  nor NOR2_561(g22536,g17076,g21911);
  nor NOR2_562(g22576,g17111,g21925);
  nor NOR2_563(g22578,g21892,g18982);
  nor NOR2_564(g22615,g21900,g18990);
  nor NOR2_565(g22651,g21912,g18997);
  nor NOR2_566(g22687,g21926,g19010);
  nor NOR2_567(g22755,g21271,g20842);
  nor NOR2_568(g22784,g16075,g20885);
  nor NOR2_569(g22789,g21278,g20850);
  nor NOR3_345(g22810,g16075,g20842,g21271);
  nor NOR2_570(g22826,g16113,g20904);
  nor NOR2_571(g22831,g21285,g20858);
  nor NOR3_346(g22851,g16113,g20850,g21278);
  nor NOR2_572(g22865,g16164,g20928);
  nor NOR2_573(g22870,g21293,g20866);
  nor NOR3_347(g22886,g16164,g20858,g21285);
  nor NOR2_574(g22900,g16223,g20956);
  nor NOR3_348(g22921,g16223,g20866,g21293);
  nor NOR2_575(g22935,g21903,g7466);
  nor NOR2_576(g22953,g20700,g7595);
  nor NOR2_577(g22985,g21618,g21049);
  nor NOR2_578(g22987,g21646,g21068);
  nor NOR2_579(g22990,g21677,g21078);
  nor NOR2_580(g22997,g21706,g21092);
  nor NOR2_581(g22999,g21085,g19241);
  nor NOR2_582(g23000,g16909,g21067);
  nor NOR2_583(g23009,g21738,g21107);
  nor NOR2_584(g23013,g21097,g19254);
  nor NOR2_585(g23014,g16939,g21077);
  nor NOR2_586(g23022,g16968,g21086);
  nor NOR3_349(g23023,g14256,g14175,g21123);
  nor NOR2_587(g23025,g21762,g21124);
  nor NOR2_588(g23029,g21111,g19267);
  nor NOR2_589(g23030,g16970,g21091);
  nor NOR2_590(g23039,g16989,g21098);
  nor NOR3_350(g23040,g14378,g14290,g21142);
  nor NOR2_591(g23042,g21778,g21143);
  nor NOR2_592(g23046,g21128,g19282);
  nor NOR2_593(g23047,g16991,g21103);
  nor NOR2_594(g23051,g21121,g21153);
  nor NOR2_595(g23058,g16999,g21112);
  nor NOR3_351(g23059,g14490,g14412,g21162);
  nor NOR2_596(g23061,g21793,g21163);
  nor NOR3_352(g23066,g21138,g19303,g19320);
  nor NOR2_597(g23067,g17015,g21122);
  nor NOR2_598(g23070,g21140,g21173);
  nor NOR2_599(g23076,g17023,g21129);
  nor NOR3_353(g23077,g14577,g14524,g21182);
  nor NOR3_354(g23080,g21158,g19324,g19347);
  nor NOR2_600(g23081,g17045,g21141);
  nor NOR2_601(g23083,g21160,g21193);
  nor NOR2_602(g23092,g17055,g21154);
  nor NOR2_603(g23093,g17056,g21155);
  nor NOR3_355(g23096,g21178,g19351,g19381);
  nor NOR2_604(g23097,g17079,g21161);
  nor NOR2_605(g23099,g21180,g21208);
  nor NOR2_606(g23110,g17090,g21174);
  nor NOR2_607(g23111,g17091,g21175);
  nor NOR3_356(g23113,g21198,g19385,g19413);
  nor NOR2_608(g23114,g17114,g21181);
  nor NOR2_609(g23117,g17117,g21188);
  nor NOR2_610(g23123,g17128,g21194);
  nor NOR2_611(g23124,g17129,g21195);
  nor NOR2_612(g23126,g17144,g21203);
  nor NOR2_613(g23132,g17155,g21209);
  nor NOR2_614(g23133,g17156,g21210);
  nor NOR2_615(g23135,g21229,g19449);
  nor NOR2_616(g23136,g20878,g10024);
  nor NOR2_617(g23137,g17167,g21218);
  nor NOR2_618(g23324,g22144,g10024);
  nor NOR2_619(g23329,g22165,g10133);
  nor NOR2_620(g23330,g22186,g22777);
  nor NOR2_621(g23339,g22181,g10238);
  nor NOR2_622(g23348,g22195,g10340);
  nor NOR2_623(g23357,g22210,g20127);
  nor NOR2_624(g23358,g22227,g18407);
  nor NOR2_625(g23359,g22216,g22907);
  nor NOR2_626(g23385,g17393,g22517);
  nor NOR2_627(g23386,g22483,g21388);
  nor NOR2_628(g23392,g17460,g22557);
  nor NOR2_629(g23393,g22526,g21418);
  nor NOR2_630(g23399,g17506,g22581);
  nor NOR2_631(g23400,g17540,g22597);
  nor NOR2_632(g23401,g22566,g21452);
  nor NOR2_633(g23406,g17597,g22618);
  nor NOR2_634(g23407,g17630,g22634);
  nor NOR2_635(g23408,g22606,g21494);
  nor NOR2_636(g23413,g17694,g22654);
  nor NOR2_637(g23418,g17794,g22690);
  nor NOR2_638(g23427,g22699,g21589);
  nor NOR2_639(g23433,g22726,g21611);
  nor NOR2_640(g23461,g22841,g21707);
  nor NOR2_641(g23477,g22906,g21758);
  nor NOR2_642(g23497,g22876,g5606);
  nor NOR2_643(g23513,g22911,g5631);
  nor NOR2_644(g23528,g22936,g5659);
  nor NOR2_645(g23539,g22942,g5697);
  nor NOR2_646(g23545,g22984,g20285);
  nor NOR3_357(g23823,g23009,g18490,g4456);
  nor NOR3_358(g23858,g23025,g18554,g4632);
  nor NOR3_359(g23892,g23042,g18604,g4809);
  nor NOR3_360(g23913,g23061,g18636,g4985);
  nor NOR2_647(g23922,g4456,g22985);
  nor NOR3_361(g23945,g4456,g13565,g23009);
  nor NOR2_648(g23950,g22992,g6707);
  nor NOR2_649(g23954,g4632,g22987);
  nor NOR3_362(g23974,g4632,g13573,g23025);
  nor NOR2_650(g23979,g23003,g7009);
  nor NOR2_651(g23983,g4809,g22990);
  nor NOR3_363(g24004,g4809,g13582,g23042);
  nor NOR2_652(g24009,g23017,g7259);
  nor NOR2_653(g24013,g4985,g22997);
  nor NOR3_364(g24038,g4985,g13602,g23061);
  nor NOR2_654(g24043,g23033,g7455);
  nor NOR2_655(g24059,g21990,g20809);
  nor NOR2_656(g24072,g22004,g20826);
  nor NOR2_657(g24083,g22015,g20836);
  nor NOR2_658(g24092,g22020,g20840);
  nor NOR2_659(g24174,g16894,g22206);
  nor NOR2_660(g24178,g16908,g22211);
  nor NOR2_661(g24179,g16923,g22214);
  nor NOR2_662(g24181,g16938,g22220);
  nor NOR2_663(g24182,g16953,g22223);
  nor NOR2_664(g24206,g16966,g22228);
  nor NOR2_665(g24207,g16967,g22229);
  nor NOR2_666(g24208,g16969,g22235);
  nor NOR2_667(g24209,g16984,g22238);
  nor NOR2_668(g24212,g16987,g22244);
  nor NOR2_669(g24213,g16988,g22245);
  nor NOR2_670(g24214,g16990,g22250);
  nor NOR2_671(g24215,g16993,g22254);
  nor NOR2_672(g24216,g16994,g22255);
  nor NOR2_673(g24218,g16997,g22264);
  nor NOR2_674(g24219,g16998,g22265);
  nor NOR2_675(g24222,g17017,g22272);
  nor NOR2_676(g24223,g17018,g22273);
  nor NOR2_677(g24225,g17021,g22281);
  nor NOR2_678(g24226,g17022,g22282);
  nor NOR2_679(g24227,g22270,g21137);
  nor NOR2_680(g24228,g17028,g22285);
  nor NOR2_681(g24230,g17047,g22291);
  nor NOR2_682(g24231,g17048,g22292);
  nor NOR2_683(g24232,g22637,g22665);
  nor NOR2_684(g24234,g22289,g21157);
  nor NOR2_685(g24235,g17062,g22305);
  nor NOR2_686(g24237,g17081,g22311);
  nor NOR2_687(g24238,g17082,g22312);
  nor NOR2_688(g24242,g22309,g21177);
  nor NOR2_689(g24243,g17097,g22333);
  nor NOR2_690(g24249,g22337,g21197);
  nor NOR2_691(g24250,g17135,g22358);
  nor NOR2_692(g24426,g23386,g10024);
  nor NOR2_693(g24428,g23544,g22398);
  nor NOR2_694(g24430,g23393,g10133);
  nor NOR2_695(g24434,g23401,g10238);
  nor NOR2_696(g24438,g23408,g10340);
  nor NOR2_697(g24445,g23427,g22777);
  nor NOR2_698(g24446,g23433,g22907);
  nor NOR2_699(g24473,g23461,g18407);
  nor NOR2_700(g24476,g23477,g20127);
  nor NOR2_701(g24479,g23593,g22516);
  nor NOR2_702(g24480,g23617,g23659);
  nor NOR2_703(g24481,g23618,g19696);
  nor NOR2_704(g24485,g23625,g22556);
  nor NOR2_705(g24486,g23643,g22577);
  nor NOR2_706(g24487,g23666,g23709);
  nor NOR2_707(g24488,g23667,g19740);
  nor NOR2_708(g24489,g23674,g22596);
  nor NOR2_709(g24490,g23686,g22607);
  nor NOR2_710(g24491,g15247,g23735);
  nor NOR2_711(g24492,g23689,g22610);
  nor NOR2_712(g24493,g23693,g22614);
  nor NOR2_713(g24494,g23716,g23763);
  nor NOR2_714(g24495,g23717,g19783);
  nor NOR2_715(g24496,g23724,g22633);
  nor NOR2_716(g24497,g23734,g22638);
  nor NOR2_717(g24498,g15324,g23777);
  nor NOR2_718(g24499,g15325,g23778);
  nor NOR2_719(g24500,g23740,g22643);
  nor NOR2_720(g24501,g15339,g23790);
  nor NOR2_721(g24502,g23743,g22646);
  nor NOR2_722(g24503,g23747,g22650);
  nor NOR2_723(g24504,g23770,g23818);
  nor NOR2_724(g24505,g23771,g19825);
  nor NOR2_725(g24506,g23776,g22667);
  nor NOR2_726(g24507,g15391,g23824);
  nor NOR2_727(g24508,g15392,g23825);
  nor NOR2_728(g24509,g23789,g22674);
  nor NOR2_729(g24510,g15410,g23830);
  nor NOR2_730(g24511,g15411,g23831);
  nor NOR2_731(g24512,g23795,g22679);
  nor NOR2_732(g24513,g15425,g23843);
  nor NOR2_733(g24514,g23798,g22682);
  nor NOR2_734(g24515,g23802,g22686);
  nor NOR2_735(g24516,g23820,g22700);
  nor NOR2_736(g24517,g23822,g22701);
  nor NOR2_737(g24519,g15459,g23855);
  nor NOR2_738(g24520,g23829,g22707);
  nor NOR2_739(g24521,g15475,g23859);
  nor NOR2_740(g24522,g15476,g23860);
  nor NOR2_741(g24523,g23842,g22714);
  nor NOR2_742(g24524,g15494,g23865);
  nor NOR2_743(g24525,g15495,g23866);
  nor NOR2_744(g24526,g23848,g22719);
  nor NOR2_745(g24527,g15509,g23878);
  nor NOR2_746(g24528,g23851,g22722);
  nor NOR2_747(g24530,g23857,g22732);
  nor NOR2_748(g24532,g15545,g23889);
  nor NOR2_749(g24533,g23864,g22738);
  nor NOR2_750(g24534,g15561,g23893);
  nor NOR2_751(g24535,g15562,g23894);
  nor NOR2_752(g24536,g23877,g22745);
  nor NOR2_753(g24537,g15580,g23899);
  nor NOR2_754(g24538,g15581,g23900);
  nor NOR2_755(g24543,g23891,g22764);
  nor NOR2_756(g24545,g15623,g23910);
  nor NOR2_757(g24546,g23898,g22770);
  nor NOR2_758(g24547,g15639,g23914);
  nor NOR2_759(g24548,g15640,g23915);
  nor NOR2_760(g24555,g23912,g22798);
  nor NOR2_761(g24557,g15699,g23942);
  nor NOR2_762(g24558,g23917,g22804);
  nor NOR2_763(g24566,g23944,g22842);
  nor NOR2_764(g24575,g23972,g22874);
  nor NOR2_765(g24606,g24183,g537);
  nor NOR2_766(g24613,g23592,g22515);
  nor NOR2_767(g24622,g23616,g22546);
  nor NOR2_768(g24623,g24183,g529);
  nor NOR2_769(g24624,g23624,g22555);
  nor NOR2_770(g24636,g24183,g530);
  nor NOR2_771(g24637,g23665,g22587);
  nor NOR2_772(g24638,g23673,g22595);
  nor NOR2_773(g24652,g24183,g531);
  nor NOR2_774(g24656,g23715,g22624);
  nor NOR2_775(g24657,g23723,g22632);
  nor NOR2_776(g24663,g24183,g532);
  nor NOR2_777(g24675,g23769,g22660);
  nor NOR2_778(g24681,g24183,g533);
  nor NOR2_779(g24682,g23688,g24183);
  nor NOR2_780(g24694,g24183,g534);
  nor NOR2_781(g24708,g23854,g22727);
  nor NOR2_782(g24711,g24183,g536);
  nor NOR2_783(g24717,g23886,g22754);
  nor NOR2_784(g24720,g23888,g22759);
  nor NOR2_785(g24728,g23907,g22788);
  nor NOR2_786(g24731,g23909,g22793);
  nor NOR2_787(g24736,g23939,g22830);
  nor NOR2_788(g24739,g23941,g22835);
  nor NOR2_789(g24742,g23971,g22869);
  nor NOR2_790(g24756,g16089,g24211);
  nor NOR2_791(g24770,g16119,g24217);
  nor NOR2_792(g24782,g16160,g24221);
  nor NOR2_793(g24783,g16161,g24224);
  nor NOR2_794(g24800,g16211,g24229);
  nor NOR2_795(g24819,g16262,g24236);
  nor NOR2_796(g24836,g16309,g24241);
  nor NOR2_797(g24845,g16350,g24246);
  nor NOR2_798(g24847,g16356,g24247);
  nor NOR2_799(g24859,g16390,g24253);
  nor NOR2_800(g24871,g16422,g24256);
  nor NOR2_801(g25027,g24227,g17001);
  nor NOR2_802(g25042,g24234,g17031);
  nor NOR2_803(g25056,g24242,g17065);
  nor NOR2_804(g25067,g24249,g17100);
  nor NOR2_805(g25075,g13880,g23483);
  nor NOR2_806(g25076,g23409,g22187);
  nor NOR2_807(g25077,g23414,g22196);
  nor NOR2_808(g25078,g23419,g22201);
  nor NOR2_809(g25081,g23423,g22202);
  nor NOR2_810(g25082,g23428,g22207);
  nor NOR2_811(g25085,g23432,g22208);
  nor NOR2_812(g25091,g23434,g22215);
  nor NOR2_813(g25099,g23440,g22224);
  nor NOR2_814(g25125,g23510,g22340);
  nor NOR2_815(g25127,g23525,g22363);
  nor NOR2_816(g25129,g23536,g22383);
  nor NOR2_817(g25185,g24492,g10024);
  nor NOR2_818(g25189,g24502,g10133);
  nor NOR2_819(g25191,g24516,g22777);
  nor NOR2_820(g25194,g24514,g10238);
  nor NOR2_821(g25197,g24528,g10340);
  nor NOR2_822(g25199,g24558,g20127);
  nor NOR2_823(g25201,g24575,g18407);
  nor NOR2_824(g25202,g24566,g22907);
  nor NOR2_825(g25204,g24745,g23547);
  nor NOR2_826(g25206,g24746,g23550);
  nor NOR2_827(g25207,g24747,g23551);
  nor NOR2_828(g25208,g24748,g23552);
  nor NOR2_829(g25209,g24749,g23554);
  nor NOR2_830(g25211,g24750,g23558);
  nor NOR2_831(g25212,g24751,g23559);
  nor NOR2_832(g25213,g24752,g23560);
  nor NOR2_833(g25214,g24754,g23563);
  nor NOR2_834(g25215,g24755,g23564);
  nor NOR2_835(g25216,g24757,g23565);
  nor NOR2_836(g25217,g24758,g23567);
  nor NOR2_837(g25218,g24760,g23571);
  nor NOR2_838(g25219,g24761,g23572);
  nor NOR2_839(g25220,g24762,g23573);
  nor NOR2_840(g25221,g24767,g23577);
  nor NOR2_841(g25222,g24768,g23578);
  nor NOR2_842(g25223,g24769,g23579);
  nor NOR2_843(g25224,g24772,g23582);
  nor NOR2_844(g25225,g24773,g23583);
  nor NOR2_845(g25226,g24774,g23584);
  nor NOR2_846(g25227,g24775,g23586);
  nor NOR2_847(g25228,g24776,g23590);
  nor NOR2_848(g25229,g24777,g23591);
  nor NOR2_849(g25230,g24779,g23598);
  nor NOR2_850(g25231,g24780,g23599);
  nor NOR2_851(g25232,g24781,g23600);
  nor NOR2_852(g25233,g24788,g23604);
  nor NOR2_853(g25234,g24789,g23605);
  nor NOR2_854(g25235,g24790,g23606);
  nor NOR2_855(g25236,g24792,g23609);
  nor NOR2_856(g25237,g24793,g23610);
  nor NOR2_857(g25238,g24794,g23611);
  nor NOR2_858(g25239,g24796,g23615);
  nor NOR2_859(g25240,g24798,g23622);
  nor NOR2_860(g25241,g24799,g23623);
  nor NOR2_861(g25242,g24802,g23630);
  nor NOR2_862(g25243,g24803,g23631);
  nor NOR2_863(g25244,g24804,g23632);
  nor NOR2_864(g25245,g24809,g23636);
  nor NOR2_865(g25246,g24810,g23637);
  nor NOR2_866(g25247,g24811,g23638);
  nor NOR2_867(g25248,g24818,g23664);
  nor NOR2_868(g25249,g24821,g23671);
  nor NOR2_869(g25250,g24822,g23672);
  nor NOR2_870(g25251,g24824,g23679);
  nor NOR2_871(g25252,g24825,g23680);
  nor NOR2_872(g25253,g24826,g23681);
  nor NOR2_873(g25254,g24831,g23687);
  nor NOR2_874(g25255,g24838,g23714);
  nor NOR2_875(g25256,g24840,g23721);
  nor NOR2_876(g25257,g24841,g23722);
  nor NOR2_877(g25258,g24846,g23741);
  nor NOR2_878(g25259,g24853,g23768);
  nor NOR2_879(g25260,g24858,g17737);
  nor NOR2_880(g25261,g24861,g23796);
  nor NOR2_881(g25262,g24869,g17824);
  nor NOR2_882(g25263,g24874,g17838);
  nor NOR2_883(g25264,g24876,g23849);
  nor NOR2_884(g25265,g24878,g23852);
  nor NOR2_885(g25266,g24881,g17912);
  nor NOR2_886(g25267,g24884,g17936);
  nor NOR2_887(g25268,g24888,g17950);
  nor NOR2_888(g25270,g24898,g18023);
  nor NOR2_889(g25271,g24901,g18047);
  nor NOR2_890(g25272,g24905,g18061);
  nor NOR2_891(g25273,g24907,g23904);
  nor NOR2_892(g25279,g24921,g18140);
  nor NOR2_893(g25280,g24924,g18164);
  nor NOR2_894(g25288,g24938,g18256);
  nor NOR2_895(g25311,g24964,g24029);
  nor NOR2_896(g25343,g24975,g5623);
  nor NOR2_897(g25357,g24986,g5651);
  nor NOR2_898(g25372,g24997,g5689);
  nor NOR2_899(g25389,g25005,g5741);
  nor NOR2_900(g25418,g24482,g22319);
  nor NOR2_901(g25426,g24183,g24616);
  nor NOR2_902(g25429,g24482,g22319);
  nor NOR2_903(g25450,g16018,g25086);
  nor NOR2_904(g25451,g16048,g25102);
  nor NOR2_905(g25452,g16101,g25117);
  nor NOR2_906(g25523,g20842,g24429);
  nor NOR2_907(g25539,g25088,g6157);
  nor NOR2_908(g25569,g24708,g24490);
  nor NOR2_909(g25589,g20850,g24433);
  nor NOR2_910(g25605,g25096,g6184);
  nor NOR2_911(g25631,g24717,g24497);
  nor NOR2_912(g25648,g24720,g24500);
  nor NOR2_913(g25668,g20858,g24437);
  nor NOR2_914(g25684,g25106,g6216);
  nor NOR2_915(g25699,g24613,g24506);
  nor NOR2_916(g25708,g24728,g24509);
  nor NOR2_917(g25725,g24731,g24512);
  nor NOR2_918(g25745,g20866,g24440);
  nor NOR2_919(g25761,g25112,g6305);
  nor NOR2_920(g25764,g25076,g21615);
  nor NOR2_921(g25772,g24624,g24520);
  nor NOR2_922(g25781,g24736,g24523);
  nor NOR2_923(g25798,g24739,g24526);
  nor NOR2_924(g25818,g25077,g21643);
  nor NOR2_925(g25826,g24638,g24533);
  nor NOR2_926(g25835,g24742,g24536);
  nor NOR3_365(g25852,g4456,g14831,g25078);
  nor NOR2_927(g25853,g25081,g21674);
  nor NOR2_928(g25861,g24657,g24546);
  nor NOR4_16(g25870,g4456,g25078,g18429,g16075);
  nor NOR3_366(g25873,g4632,g14904,g25082);
  nor NOR2_929(g25874,g25085,g21703);
  nor NOR4_17(g25882,g4632,g25082,g18502,g16113);
  nor NOR3_367(g25885,g4809,g14985,g25091);
  nor NOR4_18(g25887,g4809,g25091,g18566,g16164);
  nor NOR3_368(g25890,g4985,g15074,g25099);
  nor NOR4_19(g25892,g4985,g25099,g18616,g16223);
  nor NOR2_930(g25932,g25125,g17001);
  nor NOR2_931(g25935,g25127,g17031);
  nor NOR2_932(g25938,g25129,g17065);
  nor NOR2_933(g25940,g24428,g17100);
  nor NOR2_934(g25941,g24529,g24540);
  nor NOR2_935(g25943,g24541,g24550);
  nor NOR2_936(g25944,g24542,g24552);
  nor NOR2_937(g25946,g24553,g24561);
  nor NOR2_938(g25947,g24554,g24563);
  nor NOR2_939(g25948,g24564,g24571);
  nor NOR2_940(g25949,g24565,g24573);
  nor NOR2_941(g25950,g24574,g24580);
  nor NOR2_942(g25962,g24591,g23496);
  nor NOR2_943(g25967,g24596,g23512);
  nor NOR2_944(g25974,g24604,g23527);
  nor NOR2_945(g25979,g24611,g23538);
  nor NOR2_946(g26025,g25392,g17193);
  nor NOR2_947(g26031,g25273,g22777);
  nor NOR2_948(g26037,g25311,g18407);
  nor NOR2_949(g26041,g25475,g24855);
  nor NOR2_950(g26042,g25505,g24867);
  nor NOR2_951(g26043,g25506,g24870);
  nor NOR2_952(g26044,g25552,g24882);
  nor NOR2_953(g26045,g25553,g24885);
  nor NOR2_954(g26046,g25618,g24899);
  nor NOR2_955(g26047,g25619,g24902);
  nor NOR2_956(g26048,g25628,g24906);
  nor NOR2_957(g26049,g25629,g24908);
  nor NOR2_958(g26050,g25697,g24922);
  nor NOR2_959(g26055,g25881,g24974);
  nor NOR2_960(g26081,g25470,g25482);
  nor NOR2_961(g26083,g25426,g22319);
  nor NOR2_962(g26084,g25487,g25513);
  nor NOR3_369(g26087,g6068,g24183,g25319);
  nor NOR2_963(g26090,g25518,g25560);
  nor NOR3_370(g26096,g6068,g24183,g25394);
  nor NOR3_371(g26099,g6068,g24183,g25313);
  nor NOR2_964(g26103,g25565,g25626);
  nor NOR3_372(g26107,g6068,g24183,g25383);
  nor NOR3_373(g26110,g6068,g24183,g25305);
  nor NOR2_965(g26113,g25426,g22319);
  nor NOR3_374(g26126,g6068,g24183,g25368);
  nor NOR3_375(g26137,g6068,g24183,g25355);
  nor NOR2_966(g26140,g24183,g25430);
  nor NOR3_376(g26145,g6068,g24183,g25347);
  nor NOR3_377(g26151,g6068,g24183,g25335);
  nor NOR3_378(g26154,g6068,g24183,g25329);
  nor NOR2_967(g26160,g25951,g16162);
  nor NOR2_968(g26168,g25953,g16212);
  nor NOR2_969(g26183,g25957,g13270);
  nor NOR2_970(g26199,g25961,g13291);
  nor NOR2_971(g26217,g25963,g13320);
  nor NOR2_972(g26240,g25968,g13340);
  nor NOR2_973(g26265,g25972,g13360);
  nor NOR2_974(g26272,g25973,g16423);
  nor NOR2_975(g26283,g25954,g24486);
  nor NOR2_976(g26295,g25977,g13385);
  nor NOR2_977(g26304,g25978,g16451);
  nor NOR2_978(g26327,g25958,g24493);
  nor NOR2_979(g26336,g25981,g13481);
  nor NOR2_980(g26374,g25964,g24503);
  nor NOR2_981(g26417,g25969,g24515);
  nor NOR2_982(g26529,g25962,g17001);
  nor NOR2_983(g26530,g25967,g17031);
  nor NOR2_984(g26531,g25974,g17065);
  nor NOR2_985(g26532,g25979,g17100);
  nor NOR2_986(g26534,g25321,g8869);
  nor NOR2_987(g26541,g13755,g25269);
  nor NOR2_988(g26545,g13790,g25277);
  nor NOR2_989(g26547,g13796,g25278);
  nor NOR2_990(g26553,g13816,g25282);
  nor NOR2_991(g26557,g13818,g25286);
  nor NOR2_992(g26559,g13824,g25287);
  nor NOR2_993(g26560,g25281,g24559);
  nor NOR2_994(g26569,g13837,g25290);
  nor NOR2_995(g26573,g13839,g25294);
  nor NOR2_996(g26575,g13845,g25295);
  nor NOR2_997(g26583,g25289,g24569);
  nor NOR2_998(g26592,g13851,g25300);
  nor NOR2_999(g26596,g13853,g25304);
  nor NOR2_1000(g26607,g25299,g24578);
  nor NOR2_1001(g26616,g13860,g25310);
  nor NOR2_1002(g26630,g25309,g24585);
  nor NOR2_1003(g26655,g25328,g17084);
  nor NOR2_1004(g26659,g25334,g17116);
  nor NOR2_1005(g26660,g25208,g10024);
  nor NOR2_1006(g26661,g25337,g17122);
  nor NOR2_1007(g26664,g25346,g17138);
  nor NOR2_1008(g26665,g25348,g17143);
  nor NOR2_1009(g26666,g25216,g10133);
  nor NOR2_1010(g26667,g25351,g17149);
  nor NOR2_1011(g26669,g25360,g17161);
  nor NOR2_1012(g26670,g25362,g17166);
  nor NOR2_1013(g26671,g25226,g10238);
  nor NOR2_1014(g26672,g25365,g17172);
  nor NOR2_1015(g26675,g25375,g17176);
  nor NOR2_1016(g26676,g25377,g17181);
  nor NOR2_1017(g26677,g25238,g10340);
  nor NOR2_1018(g26776,g26042,g10024);
  nor NOR2_1019(g26781,g26044,g10133);
  nor NOR2_1020(g26786,g26049,g22777);
  nor NOR2_1021(g26789,g26046,g10238);
  nor NOR2_1022(g26795,g26050,g10340);
  nor NOR2_1023(g26798,g26055,g18407);
  nor NOR2_1024(g26799,g26158,g25453);
  nor NOR2_1025(g26800,g26163,g25457);
  nor NOR2_1026(g26801,g26171,g25461);
  nor NOR2_1027(g26802,g26188,g25466);
  nor NOR2_1028(g26803,g15105,g26213);
  nor NOR2_1029(g26804,g15172,g26235);
  nor NOR2_1030(g26805,g15173,g26236);
  nor NOR2_1031(g26806,g15197,g26244);
  nor NOR2_1032(g26807,g15245,g26261);
  nor NOR2_1033(g26808,g15246,g26262);
  nor NOR2_1034(g26809,g15258,g26270);
  nor NOR2_1035(g26810,g15259,g26271);
  nor NOR2_1036(g26811,g15283,g26279);
  nor NOR2_1037(g26812,g15321,g26291);
  nor NOR2_1038(g26813,g15337,g26302);
  nor NOR2_1039(g26814,g15338,g26303);
  nor NOR2_1040(g26815,g15350,g26311);
  nor NOR2_1041(g26816,g15351,g26312);
  nor NOR2_1042(g26817,g15375,g26317);
  nor NOR2_1043(g26818,g15407,g26335);
  nor NOR2_1044(g26820,g15423,g26346);
  nor NOR2_1045(g26821,g15424,g26347);
  nor NOR2_1046(g26822,g15436,g26352);
  nor NOR2_1047(g26823,g15437,g26353);
  nor NOR2_1048(g26824,g15491,g26382);
  nor NOR2_1049(g26825,g15507,g26390);
  nor NOR2_1050(g26826,g15508,g26391);
  nor NOR2_1051(g26827,g15577,g26425);
  nor NOR2_1052(g26869,g26458,g5642);
  nor NOR2_1053(g26873,g25483,g26260);
  nor NOR2_1054(g26877,g26140,g22319);
  nor NOR2_1055(g26878,g26482,g5680);
  nor NOR2_1056(g26882,g25514,g26301);
  nor NOR2_1057(g26885,g26140,g22319);
  nor NOR2_1058(g26887,g26498,g5732);
  nor NOR2_1059(g26891,g25561,g26345);
  nor NOR2_1060(g26897,g26513,g5790);
  nor NOR2_1061(g26901,g25627,g26389);
  nor NOR2_1062(g26905,g26096,g22319);
  nor NOR2_1063(g26914,g26107,g22319);
  nor NOR2_1064(g26988,g24893,g26023);
  nor NOR2_1065(g26989,g26663,g21913);
  nor NOR2_1066(g27011,g24916,g26026);
  nor NOR2_1067(g27012,g26668,g21931);
  nor NOR2_1068(g27037,g24933,g26028);
  nor NOR2_1069(g27038,g26674,g20640);
  nor NOR2_1070(g27051,g4456,g26081);
  nor NOR2_1071(g27065,g24945,g26029);
  nor NOR2_1072(g27066,g26024,g20665);
  nor NOR2_1073(g27078,g4632,g26084);
  nor NOR2_1074(g27094,g4809,g26090);
  nor NOR2_1075(g27106,g4985,g26103);
  nor NOR2_1076(g27120,g26560,g17001);
  nor NOR2_1077(g27123,g26583,g17031);
  nor NOR2_1078(g27129,g26607,g17065);
  nor NOR2_1079(g27131,g26630,g17100);
  nor NOR2_1080(g27144,g23451,g26052);
  nor NOR2_1081(g27147,g23458,g26054);
  nor NOR2_1082(g27149,g23462,g26060);
  nor NOR2_1083(g27152,g23467,g26062);
  nor NOR2_1084(g27157,g23471,g26067);
  nor NOR2_1085(g27160,g23476,g26069);
  nor NOR2_1086(g27165,g23484,g26074);
  nor NOR2_1087(g27174,g23494,g26080);
  nor NOR2_1088(g27175,g26075,g25342);
  nor NOR2_1089(g27179,g26082,g25356);
  nor NOR2_1090(g27184,g26085,g25371);
  nor NOR2_1091(g27188,g26091,g25388);
  nor NOR2_1092(g27243,g26802,g10340);
  nor NOR2_1093(g27250,g26955,g26166);
  nor NOR2_1094(g27251,g26958,g26186);
  nor NOR2_1095(g27252,g26963,g26207);
  nor NOR2_1096(g27253,g26965,g26212);
  nor NOR2_1097(g27254,g26968,g26231);
  nor NOR2_1098(g27255,g26969,g26233);
  nor NOR2_1099(g27256,g26970,g26234);
  nor NOR2_1100(g27257,g26971,g26243);
  nor NOR2_1101(g27258,g26977,g26257);
  nor NOR2_1102(g27259,g26978,g26258);
  nor NOR2_1103(g27260,g26979,g26259);
  nor NOR2_1104(g27261,g26980,g26263);
  nor NOR2_1105(g27262,g26981,g26268);
  nor NOR2_1106(g27263,g26982,g26269);
  nor NOR2_1107(g27264,g26984,g26278);
  nor NOR2_1108(g27265,g26993,g26288);
  nor NOR2_1109(g27266,g26994,g26289);
  nor NOR2_1110(g27267,g26995,g26290);
  nor NOR2_1111(g27268,g26996,g26292);
  nor NOR2_1112(g27269,g26997,g26293);
  nor NOR2_1113(g27270,g26998,g26298);
  nor NOR2_1114(g27271,g26999,g26299);
  nor NOR2_1115(g27272,g27000,g26300);
  nor NOR2_1116(g27273,g27001,g26307);
  nor NOR2_1117(g27274,g27002,g26309);
  nor NOR2_1118(g27275,g27003,g26310);
  nor NOR2_1119(g27276,g27004,g26316);
  nor NOR2_1120(g27277,g27005,g26318);
  nor NOR2_1121(g27278,g27006,g26319);
  nor NOR2_1122(g27279,g27007,g26324);
  nor NOR2_1123(g27280,g27008,g26325);
  nor NOR2_1124(g27281,g27009,g26326);
  nor NOR2_1125(g27282,g27016,g26332);
  nor NOR2_1126(g27283,g27017,g26333);
  nor NOR2_1127(g27284,g27018,g26334);
  nor NOR2_1128(g27285,g27019,g26339);
  nor NOR2_1129(g27286,g27020,g26340);
  nor NOR2_1130(g27287,g27021,g26342);
  nor NOR2_1131(g27288,g27022,g26343);
  nor NOR2_1132(g27289,g27023,g26344);
  nor NOR2_1133(g27290,g27024,g26348);
  nor NOR2_1134(g27291,g27025,g26350);
  nor NOR2_1135(g27292,g27026,g26351);
  nor NOR2_1136(g27293,g27027,g26357);
  nor NOR2_1137(g27294,g27028,g26361);
  nor NOR2_1138(g27295,g27029,g26362);
  nor NOR2_1139(g27296,g27030,g26363);
  nor NOR2_1140(g27297,g27031,g26365);
  nor NOR2_1141(g27298,g27032,g26366);
  nor NOR2_1142(g27299,g27033,g26371);
  nor NOR2_1143(g27300,g27034,g26372);
  nor NOR2_1144(g27301,g27035,g26373);
  nor NOR2_1145(g27302,g27042,g26379);
  nor NOR2_1146(g27303,g27043,g26380);
  nor NOR2_1147(g27304,g27044,g26381);
  nor NOR2_1148(g27305,g27045,g26383);
  nor NOR2_1149(g27306,g27046,g26384);
  nor NOR2_1150(g27307,g27047,g26386);
  nor NOR2_1151(g27308,g27048,g26387);
  nor NOR2_1152(g27309,g27049,g26388);
  nor NOR2_1153(g27310,g27050,g26392);
  nor NOR2_1154(g27311,g27053,g26396);
  nor NOR2_1155(g27312,g27054,g26397);
  nor NOR2_1156(g27313,g27055,g26400);
  nor NOR2_1157(g27314,g27056,g26404);
  nor NOR2_1158(g27315,g27057,g26405);
  nor NOR2_1159(g27316,g27058,g26406);
  nor NOR2_1160(g27317,g27059,g26408);
  nor NOR2_1161(g27318,g27060,g26409);
  nor NOR2_1162(g27319,g27061,g26414);
  nor NOR2_1163(g27320,g27062,g26415);
  nor NOR2_1164(g27321,g27063,g26416);
  nor NOR2_1165(g27322,g27070,g26422);
  nor NOR2_1166(g27323,g27071,g26423);
  nor NOR2_1167(g27324,g27072,g26424);
  nor NOR2_1168(g27325,g27073,g26426);
  nor NOR2_1169(g27326,g27074,g26427);
  nor NOR2_1170(g27327,g27077,g26432);
  nor NOR2_1171(g27328,g27080,g26437);
  nor NOR2_1172(g27329,g27081,g26438);
  nor NOR2_1173(g27330,g27082,g26441);
  nor NOR2_1174(g27331,g27083,g26445);
  nor NOR2_1175(g27332,g27084,g26446);
  nor NOR2_1176(g27333,g27085,g26447);
  nor NOR2_1177(g27334,g27086,g26449);
  nor NOR2_1178(g27335,g27087,g26450);
  nor NOR2_1179(g27336,g27088,g26455);
  nor NOR2_1180(g27337,g27089,g26456);
  nor NOR2_1181(g27338,g27090,g26457);
  nor NOR2_1182(g27339,g27093,g26464);
  nor NOR2_1183(g27340,g27096,g26469);
  nor NOR2_1184(g27341,g27097,g26470);
  nor NOR2_1185(g27342,g27098,g26473);
  nor NOR2_1186(g27343,g27099,g26477);
  nor NOR2_1187(g27344,g27100,g26478);
  nor NOR2_1188(g27345,g27101,g26479);
  nor NOR2_1189(g27346,g27105,g26488);
  nor NOR2_1190(g27347,g27108,g26493);
  nor NOR2_1191(g27348,g27109,g26494);
  nor NOR2_1192(g27354,g27112,g26504);
  nor NOR2_1193(g27414,g26770,g25187);
  nor NOR3_379(g27415,g23104,g27181,g25128);
  nor NOR2_1194(g27435,g26777,g25193);
  nor NOR3_380(g27436,g23118,g27187,g24427);
  nor NOR2_1195(g27450,g26902,g24613);
  nor NOR2_1196(g27454,g26783,g25196);
  nor NOR3_381(g27455,g23127,g26758,g24431);
  nor NOR2_1197(g27462,g26892,g24622);
  nor NOR2_1198(g27464,g27178,g25975);
  nor NOR2_1199(g27466,g26915,g24624);
  nor NOR2_1200(g27470,g26790,g25198);
  nor NOR3_382(g27471,g23138,g26764,g24435);
  nor NOR2_1201(g27478,g26754,g24432);
  nor NOR2_1202(g27481,g27182,g25980);
  nor NOR2_1203(g27482,g26906,g24637);
  nor NOR2_1204(g27485,g26928,g24638);
  nor NOR3_383(g27492,g24958,g24633,g26771);
  nor NOR2_1205(g27496,g27185,g25178);
  nor NOR2_1206(g27501,g26763,g24436);
  nor NOR2_1207(g27504,g26918,g24656);
  nor NOR2_1208(g27507,g26941,g24657);
  nor NOR3_384(g27513,g24969,g24653,g26778);
  nor NOR2_1209(g27521,g26766,g24439);
  nor NOR2_1210(g27524,g26931,g24675);
  nor NOR2_1211(g27527,g26759,g19087);
  nor NOR2_1212(g27529,g4456,g26873);
  nor NOR2_1213(g27531,g26760,g25181);
  nor NOR2_1214(g27532,g26761,g25182);
  nor NOR3_385(g27538,g24982,g24672,g26784);
  nor NOR2_1215(g27546,g26769,g24441);
  nor NOR2_1216(g27549,g26765,g19093);
  nor NOR2_1217(g27551,g4632,g26882);
  nor NOR3_386(g27558,g24993,g24691,g26791);
  nor NOR2_1218(g27563,g26922,g24708);
  nor NOR2_1219(g27564,g26767,g25184);
  nor NOR2_1220(g27565,g26768,g19100);
  nor NOR2_1221(g27567,g4809,g26891);
  nor NOR2_1222(g27572,g26911,g24717);
  nor NOR2_1223(g27573,g26773,g25188);
  nor NOR2_1224(g27574,g26935,g24720);
  nor NOR2_1225(g27575,g26774,g19107);
  nor NOR2_1226(g27577,g4985,g26901);
  nor NOR2_1227(g27579,g26775,g25192);
  nor NOR2_1228(g27581,g26925,g24728);
  nor NOR2_1229(g27582,g26944,g24731);
  nor NOR2_1230(g27584,g26938,g24736);
  nor NOR2_1231(g27585,g26950,g24739);
  nor NOR2_1232(g27588,g26947,g24742);
  nor NOR2_1233(g27594,g27175,g17001);
  nor NOR2_1234(g27603,g27179,g17031);
  nor NOR2_1235(g27612,g27184,g17065);
  nor NOR2_1236(g27621,g27188,g17100);
  nor NOR2_1237(g27629,g26829,g26051);
  nor NOR2_1238(g27631,g26833,g26053);
  nor NOR2_1239(g27655,g26842,g26061);
  nor NOR2_1240(g27658,g26851,g26068);
  nor NOR2_1241(g27672,g26799,g10024);
  nor NOR2_1242(g27678,g26800,g10133);
  nor NOR2_1243(g27682,g26801,g10238);
  nor NOR2_1244(g27718,g27251,g10133);
  nor NOR2_1245(g27722,g27252,g10238);
  nor NOR2_1246(g27724,g27254,g10340);
  nor NOR2_1247(g27735,g27394,g26961);
  nor NOR2_1248(g27736,g27396,g26962);
  nor NOR2_1249(g27741,g27407,g26966);
  nor NOR2_1250(g27742,g27409,g26967);
  nor NOR2_1251(g27746,g27425,g26972);
  nor NOR2_1252(g27747,g27427,g26973);
  nor NOR2_1253(g27754,g27446,g26985);
  nor NOR2_1254(g27755,g27448,g26986);
  nor NOR2_1255(g27759,g27495,g27052);
  nor NOR2_1256(g27760,g27509,g27076);
  nor NOR2_1257(g27761,g27516,g27079);
  nor NOR2_1258(g27762,g27530,g27091);
  nor NOR2_1259(g27763,g27534,g27092);
  nor NOR2_1260(g27764,g27541,g27095);
  nor NOR2_1261(g27765,g27552,g27103);
  nor NOR2_1262(g27766,g27554,g27104);
  nor NOR2_1263(g27767,g27561,g27107);
  nor NOR2_1264(g27768,g27568,g27110);
  nor NOR2_1265(g27769,g27570,g27111);
  nor NOR2_1266(g27771,g27578,g27115);
  nor NOR2_1267(g27798,g27632,g1223);
  nor NOR3_387(g27802,g6087,g27632,g25330);
  nor NOR2_1268(g27810,g27632,g1215);
  nor NOR3_388(g27811,g6087,g27632,g25404);
  nor NOR3_389(g27814,g6087,g27632,g25322);
  nor NOR2_1269(g27823,g27632,g1216);
  nor NOR3_390(g27824,g6087,g27632,g25399);
  nor NOR3_391(g27827,g6087,g27632,g25314);
  nor NOR2_1270(g27834,g27478,g14630);
  nor NOR2_1271(g27842,g27632,g1217);
  nor NOR2_1272(g27850,g27501,g14650);
  nor NOR2_1273(g27854,g27632,g1218);
  nor NOR3_392(g27855,g6087,g27632,g25385);
  nor NOR2_1274(g27864,g27632,g1219);
  nor NOR3_393(g27865,g6087,g27632,g25370);
  nor NOR2_1275(g27868,g23742,g27632);
  nor NOR2_1276(g27869,g27632,g25437);
  nor NOR2_1277(g27875,g27521,g14677);
  nor NOR2_1278(g27882,g27632,g1220);
  nor NOR3_394(g27883,g6087,g27632,g25361);
  nor NOR2_1279(g27886,g27632,g24627);
  nor NOR2_1280(g27892,g27546,g14711);
  nor NOR2_1281(g27896,g27632,g1222);
  nor NOR3_395(g27897,g6087,g27632,g25349);
  nor NOR3_396(g27900,g6087,g27632,g25338);
  nor NOR2_1282(g27906,g16127,g27656);
  nor NOR2_1283(g27911,g16170,g27657);
  nor NOR2_1284(g27916,g16219,g27659);
  nor NOR2_1285(g27917,g16220,g27660);
  nor NOR2_1286(g27925,g16276,g27661);
  nor NOR2_1287(g27937,g16321,g27666);
  nor NOR2_1288(g27950,g16367,g27673);
  nor NOR2_1289(g27962,g16394,g27679);
  nor NOR2_1290(g27964,g16400,g27680);
  nor NOR2_1291(g27980,g16428,g27681);
  nor NOR2_1292(g27997,g16456,g27242);
  nor NOR2_1293(g28002,g26032,g27246);
  nor NOR2_1294(g28029,g26033,g27247);
  nor NOR2_1295(g28059,g26034,g27248);
  nor NOR2_1296(g28088,g26036,g27249);
  nor NOR2_1297(g28145,g27629,g17001);
  nor NOR2_1298(g28146,g27631,g17031);
  nor NOR2_1299(g28147,g27655,g17065);
  nor NOR2_1300(g28148,g27658,g17100);
  nor NOR2_1301(g28157,g13902,g27370);
  nor NOR2_1302(g28185,g27356,g26845);
  nor NOR2_1303(g28189,g27359,g26853);
  nor NOR2_1304(g28191,g27365,g26860);
  nor NOR2_1305(g28192,g27372,g26866);
  nor NOR2_1306(g28199,g27250,g10024);
  nor NOR2_1307(g28321,g27742,g10133);
  nor NOR2_1308(g28325,g27747,g10238);
  nor NOR2_1309(g28328,g27755,g10340);
  nor NOR2_1310(g28342,g15460,g28008);
  nor NOR2_1311(g28344,g15526,g28027);
  nor NOR2_1312(g28345,g15527,g28028);
  nor NOR2_1313(g28346,g15546,g28035);
  nor NOR2_1314(g28348,g15594,g28050);
  nor NOR2_1315(g28349,g15595,g28051);
  nor NOR2_1316(g28350,g15604,g28057);
  nor NOR2_1317(g28351,g15605,g28058);
  nor NOR2_1318(g28352,g15624,g28065);
  nor NOR2_1319(g28353,g15666,g28073);
  nor NOR2_1320(g28354,g15670,g28079);
  nor NOR2_1321(g28355,g15671,g28080);
  nor NOR2_1322(g28356,g15680,g28086);
  nor NOR2_1323(g28357,g15681,g28087);
  nor NOR2_1324(g28358,g15700,g28094);
  nor NOR2_1325(g28360,g15725,g28098);
  nor NOR2_1326(g28361,g15729,g28104);
  nor NOR2_1327(g28362,g15730,g28105);
  nor NOR2_1328(g28363,g15739,g28111);
  nor NOR2_1329(g28364,g15740,g28112);
  nor NOR2_1330(g28366,g15765,g28116);
  nor NOR2_1331(g28367,g15769,g28122);
  nor NOR2_1332(g28368,g15770,g28123);
  nor NOR2_1333(g28371,g15793,g28127);
  nor NOR2_1334(g28392,g27886,g22344);
  nor NOR2_1335(g28394,g27869,g22344);
  nor NOR2_1336(g28397,g27869,g22344);
  nor NOR2_1337(g28400,g27886,g22344);
  nor NOR2_1338(g28403,g27811,g22344);
  nor NOR2_1339(g28406,g27824,g22344);
  nor NOR2_1340(g28409,g24676,g27801);
  nor NOR2_1341(g28410,g27748,g22344);
  nor NOR2_1342(g28413,g24695,g27809);
  nor NOR2_1343(g28414,g27748,g22344);
  nor NOR2_1344(g28417,g24712,g27830);
  nor NOR2_1345(g28418,g24723,g27846);
  nor NOR2_1346(g28420,g16031,g28171);
  nor NOR2_1347(g28421,g16068,g28176);
  nor NOR2_1348(g28425,g16133,g28188);
  nor NOR2_1349(g28449,g27727,g26780);
  nor NOR2_1350(g28461,g27729,g26787);
  nor NOR2_1351(g28470,g27671,g28193);
  nor NOR2_1352(g28473,g27730,g26794);
  nor NOR2_1353(g28482,g27731,g26797);
  nor NOR2_1354(g28488,g26755,g27719);
  nor NOR2_1355(g28489,g26756,g27720);
  nor NOR2_1356(g28490,g27240,g27721);
  nor NOR2_1357(g28495,g27244,g27723);
  nor NOR2_1358(g28499,g26027,g27725);
  nor NOR2_1359(g28523,g26035,g27732);
  nor NOR2_1360(g28525,g27245,g27726);
  nor NOR2_1361(g28528,g26030,g27728);
  nor NOR2_1362(g28551,g26038,g27733);
  nor NOR2_1363(g28578,g26039,g27734);
  nor NOR2_1364(g28606,g26040,g27737);
  nor NOR2_1365(g28634,g28185,g17001);
  nor NOR2_1366(g28635,g28189,g17031);
  nor NOR2_1367(g28636,g28191,g17065);
  nor NOR2_1368(g28637,g28192,g17100);
  nor NOR2_1369(g28654,g27770,g27355);
  nor NOR2_1370(g28656,g27772,g27358);
  nor NOR2_1371(g28658,g27773,g27364);
  nor NOR2_1372(g28661,g27775,g27371);
  nor NOR2_1373(g28668,g27736,g10024);
  nor NOR2_1374(g28728,g28422,g27904);
  nor NOR2_1375(g28731,g28423,g27908);
  nor NOR2_1376(g28732,g14894,g28426);
  nor NOR2_1377(g28733,g28424,g27909);
  nor NOR2_1378(g28735,g14957,g28430);
  nor NOR2_1379(g28736,g28427,g27913);
  nor NOR2_1380(g28737,g28428,g27914);
  nor NOR2_1381(g28738,g14975,g28433);
  nor NOR2_1382(g28739,g28429,g27915);
  nor NOR2_1383(g28744,g15030,g28439);
  nor NOR2_1384(g28745,g28431,g27922);
  nor NOR2_1385(g28746,g15046,g28441);
  nor NOR2_1386(g28747,g28434,g27923);
  nor NOR2_1387(g28748,g28435,g27924);
  nor NOR2_1388(g28749,g15064,g28444);
  nor NOR2_1389(g28750,g28436,g27926);
  nor NOR2_1390(g28754,g28440,g27931);
  nor NOR2_1391(g28758,g15126,g28451);
  nor NOR2_1392(g28759,g28442,g27935);
  nor NOR2_1393(g28760,g15142,g28453);
  nor NOR2_1394(g28761,g28445,g27936);
  nor NOR2_1395(g28762,g28446,g27938);
  nor NOR2_1396(g28763,g15160,g28456);
  nor NOR2_1397(g28767,g28452,g27945);
  nor NOR2_1398(g28771,g15218,g28463);
  nor NOR2_1399(g28772,g28454,g27949);
  nor NOR2_1400(g28773,g15234,g28465);
  nor NOR2_1401(g28774,g28457,g27951);
  nor NOR2_1402(g28778,g28464,g27963);
  nor NOR2_1403(g28782,g15304,g28475);
  nor NOR2_1404(g28783,g28466,g27968);
  nor NOR2_1405(g28784,g28468,g27970);
  nor NOR2_1406(g28788,g28476,g27984);
  nor NOR2_1407(g28789,g28477,g27985);
  nor NOR2_1408(g28790,g28478,g27991);
  nor NOR2_1409(g28794,g28484,g28009);
  nor NOR2_1410(g28795,g28485,g28015);
  nor NOR2_1411(g28802,g28492,g28036);
  nor NOR2_1412(g28803,g28493,g28042);
  nor NOR2_1413(g28813,g28497,g28066);
  nor NOR2_1414(g28874,g28657,g16221);
  nor NOR2_1415(g28886,g28659,g16277);
  nor NOR2_1416(g28903,g28660,g13295);
  nor NOR2_1417(g28920,g28662,g13322);
  nor NOR2_1418(g28941,g28663,g13343);
  nor NOR3_397(g28954,g26673,g27241,g28323);
  nor NOR2_1419(g28963,g28664,g13365);
  nor NOR2_1420(g28982,g28665,g28670);
  nor NOR2_1421(g28987,g28666,g13390);
  nor NOR2_1422(g28990,g28667,g16457);
  nor NOR2_1423(g29009,g28669,g28320);
  nor NOR2_1424(g29013,g28671,g11607);
  nor NOR2_1425(g29016,g28672,g13487);
  nor NOR2_1426(g29031,g28319,g28324);
  nor NOR2_1427(g29039,g28322,g13500);
  nor NOR2_1428(g29063,g28326,g28329);
  nor NOR2_1429(g29064,g28327,g28330);
  nor NOR2_1430(g29083,g28331,g28333);
  nor NOR2_1431(g29090,g28332,g28334);
  nor NOR2_1432(g29097,g28335,g28336);
  nor NOR2_1433(g29109,g28654,g17001);
  nor NOR2_1434(g29110,g28656,g17031);
  nor NOR2_1435(g29111,g28658,g17065);
  nor NOR2_1436(g29112,g28661,g17100);
  nor NOR2_1437(g29113,g28381,g8907);
  nor NOR2_1438(g29126,g28373,g27774);
  nor NOR2_1439(g29127,g28376,g27779);
  nor NOR2_1440(g29128,g28380,g27783);
  nor NOR2_1441(g29129,g28385,g27790);
  nor NOR2_1442(g29167,g28841,g28396);
  nor NOR2_1443(g29169,g28843,g28398);
  nor NOR2_1444(g29170,g28844,g28399);
  nor NOR2_1445(g29172,g28846,g28401);
  nor NOR2_1446(g29173,g28847,g28402);
  nor NOR2_1447(g29178,g28848,g28404);
  nor NOR2_1448(g29179,g28849,g28405);
  nor NOR2_1449(g29181,g28850,g28407);
  nor NOR2_1450(g29182,g28851,g28408);
  nor NOR2_1451(g29184,g28852,g28411);
  nor NOR2_1452(g29185,g28853,g28412);
  nor NOR2_1453(g29187,g28854,g28416);
  nor NOR2_1454(g29194,g14958,g28881);
  nor NOR2_1455(g29195,g28880,g28438);
  nor NOR2_1456(g29197,g15031,g28893);
  nor NOR2_1457(g29198,g15047,g28898);
  nor NOR2_1458(g29199,g28892,g28448);
  nor NOR2_1459(g29201,g15104,g28910);
  nor NOR2_1460(g29202,g28897,g28450);
  nor NOR2_1461(g29204,g15127,g28915);
  nor NOR2_1462(g29205,g15143,g28923);
  nor NOR2_1463(g29206,g28909,g28459);
  nor NOR2_1464(g29207,g28914,g28460);
  nor NOR2_1465(g29209,g15196,g28936);
  nor NOR2_1466(g29210,g28919,g28462);
  nor NOR2_1467(g29212,g15219,g28944);
  nor NOR2_1468(g29213,g15235,g28949);
  nor NOR2_1469(g29214,g28931,g28469);
  nor NOR2_1470(g29215,g28935,g28471);
  nor NOR2_1471(g29216,g28940,g28472);
  nor NOR2_1472(g29218,g15282,g28966);
  nor NOR2_1473(g29219,g28948,g28474);
  nor NOR2_1474(g29221,g15305,g28971);
  nor NOR2_1475(g29222,g28958,g28479);
  nor NOR2_1476(g29223,g28962,g28480);
  nor NOR2_1477(g29224,g28970,g28481);
  nor NOR2_1478(g29226,g15374,g28997);
  nor NOR2_1479(g29227,g28986,g28486);
  nor NOR2_1480(g29228,g28996,g28487);
  nor NOR2_1481(g29231,g29022,g28494);
  nor NOR2_1482(g29303,g28716,g19112);
  nor NOR2_1483(g29313,g28717,g19117);
  nor NOR2_1484(g29324,g28718,g19124);
  nor NOR2_1485(g29333,g28719,g19131);
  nor NOR2_1486(g29340,g28337,g28722);
  nor NOR2_1487(g29343,g28338,g28724);
  nor NOR2_1488(g29345,g28339,g28726);
  nor NOR2_1489(g29347,g28340,g28729);
  nor NOR2_1490(g29353,g29126,g17001);
  nor NOR2_1491(g29354,g29127,g17031);
  nor NOR2_1492(g29355,g29128,g17065);
  nor NOR2_1493(g29357,g29129,g17100);
  nor NOR2_1494(g29399,g28834,g28378);
  nor NOR2_1495(g29403,g28836,g28383);
  nor NOR2_1496(g29406,g28838,g28387);
  nor NOR2_1497(g29409,g28840,g28389);
  nor NOR2_1498(g29552,g29130,g29411);
  nor NOR2_1499(g29569,g28708,g29174);
  nor NOR2_1500(g29570,g28709,g29175);
  nor NOR2_1501(g29571,g28710,g29176);
  nor NOR2_1502(g29574,g28712,g29180);
  nor NOR2_1503(g29576,g28713,g29183);
  nor NOR2_1504(g29577,g28714,g29186);
  nor NOR2_1505(g29578,g28715,g29188);
  nor NOR2_1506(g29579,g29399,g17001);
  nor NOR2_1507(g29580,g29403,g17031);
  nor NOR2_1508(g29581,g29406,g17065);
  nor NOR2_1509(g29582,g29409,g17100);
  nor NOR2_1510(g29606,g13878,g29248);
  nor NOR2_1511(g29608,g13892,g29251);
  nor NOR2_1512(g29609,g13900,g29252);
  nor NOR2_1513(g29611,g13913,g29255);
  nor NOR2_1514(g29612,g13933,g29256);
  nor NOR2_1515(g29613,g13941,g29257);
  nor NOR2_1516(g29616,g13969,g29259);
  nor NOR2_1517(g29617,g13989,g29260);
  nor NOR2_1518(g29618,g13997,g29261);
  nor NOR2_1519(g29620,g14039,g29262);
  nor NOR2_1520(g29621,g14059,g29263);
  nor NOR2_1521(g29623,g14130,g29264);
  nor NOR2_1522(g29663,g29518,g29284);
  nor NOR2_1523(g29665,g29521,g29289);
  nor NOR2_1524(g29667,g29524,g29294);
  nor NOR2_1525(g29669,g29528,g29300);
  nor NOR2_1526(g29670,g29529,g29302);
  nor NOR2_1527(g29671,g29534,g29310);
  nor NOR2_1528(g29672,g29536,g29312);
  nor NOR2_1529(g29676,g29540,g29320);
  nor NOR2_1530(g29677,g29543,g29321);
  nor NOR2_1531(g29678,g29545,g29323);
  nor NOR2_1532(g29679,g29549,g29329);
  nor NOR2_1533(g29680,g29553,g29330);
  nor NOR2_1534(g29681,g29555,g29332);
  nor NOR2_1535(g29682,g29557,g29336);
  nor NOR2_1536(g29683,g29559,g29337);
  nor NOR2_1537(g29684,g29562,g29338);
  nor NOR2_1538(g29685,g29564,g29341);
  nor NOR2_1539(g29686,g29566,g29342);
  nor NOR2_1540(g29687,g29572,g29344);
  nor NOR2_1541(g29688,g29575,g29346);
  nor NOR2_1542(g29703,g29583,g1917);
  nor NOR3_398(g29705,g6104,g29583,g25339);
  nor NOR2_1543(g29709,g29583,g1909);
  nor NOR3_399(g29710,g6104,g29583,g25412);
  nor NOR3_400(g29713,g6104,g29583,g25332);
  nor NOR2_1544(g29717,g29583,g1910);
  nor NOR3_401(g29718,g6104,g29583,g25409);
  nor NOR3_402(g29721,g6104,g29583,g25323);
  nor NOR2_1545(g29725,g29583,g1911);
  nor NOR2_1546(g29727,g29583,g1912);
  nor NOR3_403(g29728,g6104,g29583,g25401);
  nor NOR2_1547(g29731,g29583,g1913);
  nor NOR3_404(g29732,g6104,g29583,g25387);
  nor NOR2_1548(g29735,g23797,g29583);
  nor NOR2_1549(g29736,g29583,g25444);
  nor NOR2_1550(g29740,g29583,g1914);
  nor NOR3_405(g29741,g6104,g29583,g25376);
  nor NOR2_1551(g29744,g29583,g24641);
  nor NOR2_1552(g29747,g29583,g1916);
  nor NOR3_406(g29748,g6104,g29583,g25363);
  nor NOR3_407(g29751,g6104,g29583,g25352);
  nor NOR2_1553(g29754,g16178,g29607);
  nor NOR2_1554(g29755,g16229,g29610);
  nor NOR2_1555(g29756,g16284,g29614);
  nor NOR2_1556(g29757,g16285,g29615);
  nor NOR2_1557(g29758,g16335,g29619);
  nor NOR2_1558(g29759,g16379,g29622);
  nor NOR2_1559(g29760,g16411,g29624);
  nor NOR3_408(g29761,g28707,g28711,g29466);
  nor NOR2_1560(g29762,g16432,g29625);
  nor NOR2_1561(g29763,g16438,g29626);
  nor NOR2_1562(g29764,g16462,g29464);
  nor NOR2_1563(g29765,g13492,g29465);
  nor NOR2_1564(g29766,g29467,g19142);
  nor NOR2_1565(g29767,g29468,g19143);
  nor NOR2_1566(g29768,g29469,g19146);
  nor NOR2_1567(g29769,g29470,g19148);
  nor NOR2_1568(g29770,g29471,g29196);
  nor NOR2_1569(g29771,g29472,g29200);
  nor NOR2_1570(g29772,g29473,g29203);
  nor NOR2_1571(g29773,g29474,g29208);
  nor NOR2_1572(g29774,g29475,g29211);
  nor NOR2_1573(g29775,g29476,g29217);
  nor NOR2_1574(g29776,g29477,g29220);
  nor NOR2_1575(g29777,g29478,g29225);
  nor NOR2_1576(g29778,g29479,g29229);
  nor NOR2_1577(g29779,g13943,g29502);
  nor NOR2_1578(g29780,g29480,g29232);
  nor NOR2_1579(g29781,g29481,g29233);
  nor NOR2_1580(g29782,g29482,g29234);
  nor NOR2_1581(g29783,g29483,g29235);
  nor NOR2_1582(g29784,g29484,g29236);
  nor NOR2_1583(g29785,g29485,g29238);
  nor NOR2_1584(g29786,g29486,g29239);
  nor NOR2_1585(g29787,g29487,g29240);
  nor NOR2_1586(g29788,g29488,g29241);
  nor NOR2_1587(g29789,g29489,g29242);
  nor NOR2_1588(g29791,g29490,g29243);
  nor NOR2_1589(g29912,g24676,g29716);
  nor NOR2_1590(g29914,g24695,g29724);
  nor NOR2_1591(g29916,g24712,g29726);
  nor NOR2_1592(g29918,g29744,g22367);
  nor NOR2_1593(g29919,g29736,g22367);
  nor NOR2_1594(g29920,g24723,g29739);
  nor NOR2_1595(g29921,g29736,g22367);
  nor NOR2_1596(g29922,g29744,g22367);
  nor NOR2_1597(g29924,g29710,g22367);
  nor NOR2_1598(g29926,g29718,g22367);
  nor NOR2_1599(g29928,g29673,g22367);
  nor NOR2_1600(g29929,g29673,g22367);
  nor NOR2_1601(g29936,g16049,g29790);
  nor NOR2_1602(g29939,g16102,g29792);
  nor NOR2_1603(g29941,g16182,g29793);
  nor NOR2_1604(g30010,g29520,g29942);
  nor NOR2_1605(g30011,g29522,g29944);
  nor NOR2_1606(g30012,g29523,g29945);
  nor NOR2_1607(g30013,g29525,g29946);
  nor NOR2_1608(g30014,g29526,g29947);
  nor NOR2_1609(g30015,g29527,g29948);
  nor NOR2_1610(g30016,g29531,g29949);
  nor NOR2_1611(g30017,g29532,g29950);
  nor NOR2_1612(g30018,g29533,g29951);
  nor NOR2_1613(g30019,g29538,g29952);
  nor NOR2_1614(g30020,g29539,g29953);
  nor NOR2_1615(g30021,g29541,g29954);
  nor NOR2_1616(g30022,g29547,g29955);
  nor NOR2_1617(g30023,g29548,g29956);
  nor NOR2_1618(g30024,g29550,g29957);
  nor NOR2_1619(g30025,g29558,g29958);
  nor NOR2_1620(g30026,g29560,g29959);
  nor NOR2_1621(g30027,g29565,g29960);
  nor NOR2_1622(g30028,g29567,g29961);
  nor NOR2_1623(g30029,g29573,g29962);
  nor NOR2_1624(g30030,g24676,g29923);
  nor NOR2_1625(g30031,g24695,g29925);
  nor NOR2_1626(g30032,g24712,g29927);
  nor NOR2_1627(g30033,g24723,g29931);
  nor NOR2_1628(g30053,g29963,g16286);
  nor NOR2_1629(g30054,g29964,g16336);
  nor NOR2_1630(g30055,g29965,g13326);
  nor NOR2_1631(g30056,g29966,g13345);
  nor NOR2_1632(g30057,g29967,g13368);
  nor NOR2_1633(g30058,g29968,g13395);
  nor NOR2_1634(g30059,g29969,g29811);
  nor NOR2_1635(g30060,g29970,g11612);
  nor NOR2_1636(g30061,g29971,g13493);
  nor NOR2_1637(g30062,g29810,g29815);
  nor NOR2_1638(g30063,g29812,g11637);
  nor NOR2_1639(g30064,g29813,g13506);
  nor NOR2_1640(g30065,g29814,g29817);
  nor NOR2_1641(g30066,g29816,g13517);
  nor NOR2_1642(g30067,g29818,g29820);
  nor NOR2_1643(g30068,g29819,g29821);
  nor NOR2_1644(g30069,g29822,g29828);
  nor NOR2_1645(g30070,g29827,g29833);
  nor NOR2_1646(g30071,g29834,g29839);
  nor NOR2_1647(g30072,g29910,g8947);
  nor NOR2_1648(g30245,g16074,g30077);
  nor NOR2_1649(g30246,g16107,g30079);
  nor NOR2_1650(g30247,g16112,g30080);
  nor NOR2_1651(g30248,g16139,g30081);
  nor NOR2_1652(g30249,g16158,g30082);
  nor NOR2_1653(g30250,g16163,g30083);
  nor NOR2_1654(g30251,g16198,g30085);
  nor NOR2_1655(g30252,g16217,g30086);
  nor NOR2_1656(g30253,g16222,g30087);
  nor NOR2_1657(g30254,g16242,g30088);
  nor NOR2_1658(g30255,g16263,g30089);
  nor NOR2_1659(g30256,g16282,g30090);
  nor NOR2_1660(g30257,g16290,g30091);
  nor NOR2_1661(g30258,g16291,g30092);
  nor NOR2_1662(g30259,g16301,g30093);
  nor NOR2_1663(g30260,g16322,g30094);
  nor NOR2_1664(g30261,g16342,g30095);
  nor NOR2_1665(g30262,g16343,g30096);
  nor NOR2_1666(g30263,g16344,g30097);
  nor NOR2_1667(g30264,g16348,g30098);
  nor NOR2_1668(g30265,g16349,g30099);
  nor NOR2_1669(g30266,g16359,g30100);
  nor NOR2_1670(g30267,g16380,g30101);
  nor NOR2_1671(g30268,g16382,g30102);
  nor NOR2_1672(g30269,g16386,g30103);
  nor NOR2_1673(g30270,g16387,g30104);
  nor NOR2_1674(g30271,g16388,g30105);
  nor NOR2_1675(g30272,g16392,g30106);
  nor NOR2_1676(g30273,g16393,g30107);
  nor NOR2_1677(g30274,g16403,g30108);
  nor NOR2_1678(g30275,g16413,g30109);
  nor NOR2_1679(g30276,g16415,g30110);
  nor NOR2_1680(g30277,g16418,g30111);
  nor NOR2_1681(g30278,g16420,g30112);
  nor NOR2_1682(g30279,g16424,g30113);
  nor NOR2_1683(g30280,g16425,g30114);
  nor NOR2_1684(g30281,g16426,g30115);
  nor NOR2_1685(g30282,g16430,g30117);
  nor NOR2_1686(g30283,g16431,g30118);
  nor NOR2_1687(g30284,g16444,g29980);
  nor NOR2_1688(g30285,g16447,g29981);
  nor NOR2_1689(g30286,g16449,g29982);
  nor NOR2_1690(g30287,g16452,g29983);
  nor NOR2_1691(g30288,g16454,g29984);
  nor NOR2_1692(g30289,g16458,g29985);
  nor NOR2_1693(g30290,g16459,g29986);
  nor NOR2_1694(g30291,g16460,g29987);
  nor NOR2_1695(g30292,g13477,g29988);
  nor NOR2_1696(g30293,g13480,g29989);
  nor NOR2_1697(g30294,g13483,g29990);
  nor NOR2_1698(g30295,g13485,g29991);
  nor NOR2_1699(g30296,g13488,g29993);
  nor NOR2_1700(g30297,g13490,g29994);
  nor NOR2_1701(g30298,g13496,g29995);
  nor NOR2_1702(g30299,g13499,g29996);
  nor NOR2_1703(g30300,g13502,g30001);
  nor NOR2_1704(g30301,g13504,g30002);
  nor NOR2_1705(g30302,g13513,g30003);
  nor NOR2_1706(g30303,g13516,g30005);
  nor NOR2_1707(g30304,g13527,g30007);
  nor NOR2_1708(g30338,g14297,g30225);
  nor NOR2_1709(g30341,g14328,g30226);
  nor NOR2_1710(g30356,g14419,g30227);
  nor NOR2_1711(g30399,g30116,g30123);
  nor NOR2_1712(g30400,g29997,g30127);
  nor NOR2_1713(g30401,g29998,g30128);
  nor NOR2_1714(g30402,g29999,g30129);
  nor NOR2_1715(g30403,g30004,g30131);
  nor NOR2_1716(g30404,g30006,g30132);
  nor NOR2_1717(g30405,g30008,g30133);
  nor NOR2_1718(g30406,g30009,g30138);
  nor NOR2_1719(g30455,g13953,g30216);
  nor NOR2_1720(g30468,g14007,g30217);
  nor NOR2_1721(g30470,g14023,g30218);
  nor NOR2_1722(g30482,g14067,g30219);
  nor NOR2_1723(g30485,g14098,g30220);
  nor NOR2_1724(g30487,g14114,g30221);
  nor NOR2_1725(g30500,g14182,g30222);
  nor NOR2_1726(g30503,g14213,g30223);
  nor NOR2_1727(g30505,g14229,g30224);
  nor NOR2_1728(g30566,g14327,g30398);
  nor NOR2_1729(g30584,g30412,g2611);
  nor NOR3_409(g30588,g6119,g30412,g25353);
  nor NOR2_1730(g30593,g30412,g2603);
  nor NOR3_410(g30594,g6119,g30412,g25419);
  nor NOR3_411(g30597,g6119,g30412,g25341);
  nor NOR2_1731(g30601,g30412,g2604);
  nor NOR3_412(g30602,g6119,g30412,g25417);
  nor NOR3_413(g30605,g6119,g30412,g25333);
  nor NOR2_1732(g30608,g30412,g2605);
  nor NOR2_1733(g30609,g30412,g2606);
  nor NOR3_414(g30610,g6119,g30412,g25411);
  nor NOR2_1734(g30613,g30412,g2607);
  nor NOR3_415(g30614,g6119,g30412,g25403);
  nor NOR2_1735(g30617,g23850,g30412);
  nor NOR2_1736(g30618,g30412,g25449);
  nor NOR2_1737(g30621,g30412,g2608);
  nor NOR3_416(g30622,g6119,g30412,g25393);
  nor NOR2_1738(g30625,g30412,g24660);
  nor NOR2_1739(g30628,g30412,g2610);
  nor NOR3_417(g30629,g6119,g30412,g25378);
  nor NOR3_418(g30632,g6119,g30412,g25366);
  nor NOR2_1740(g30635,g16108,g30407);
  nor NOR2_1741(g30636,g16140,g30409);
  nor NOR2_1742(g30637,g16141,g30410);
  nor NOR2_1743(g30638,g16159,g30411);
  nor NOR2_1744(g30639,g16186,g30436);
  nor NOR2_1745(g30640,g16187,g30437);
  nor NOR2_1746(g30641,g16188,g30438);
  nor NOR2_1747(g30642,g16199,g30440);
  nor NOR2_1748(g30643,g16200,g30441);
  nor NOR2_1749(g30644,g16218,g30442);
  nor NOR2_1750(g30645,g16240,g30444);
  nor NOR2_1751(g30646,g16241,g30445);
  nor NOR2_1752(g30647,g16251,g30447);
  nor NOR2_1753(g30648,g16252,g30448);
  nor NOR2_1754(g30649,g16253,g30449);
  nor NOR2_1755(g30650,g16264,g30451);
  nor NOR2_1756(g30651,g16265,g30452);
  nor NOR2_1757(g30652,g16283,g30453);
  nor NOR2_1758(g30653,g16289,g30454);
  nor NOR2_1759(g30654,g16299,g30457);
  nor NOR2_1760(g30655,g16300,g30458);
  nor NOR2_1761(g30656,g16310,g30460);
  nor NOR2_1762(g30657,g16311,g30461);
  nor NOR2_1763(g30658,g16312,g30462);
  nor NOR2_1764(g30659,g16323,g30464);
  nor NOR2_1765(g30660,g16324,g30465);
  nor NOR2_1766(g30661,g16345,g30467);
  nor NOR2_1767(g30662,g16347,g30469);
  nor NOR2_1768(g30663,g16357,g30472);
  nor NOR2_1769(g30664,g16358,g30473);
  nor NOR2_1770(g30665,g16368,g30475);
  nor NOR2_1771(g30666,g16369,g30476);
  nor NOR2_1772(g30667,g16370,g30477);
  nor NOR2_1773(g30668,g16381,g30478);
  nor NOR2_1774(g30669,g16383,g30481);
  nor NOR2_1775(g30670,g16389,g30484);
  nor NOR2_1776(g30671,g16391,g30486);
  nor NOR2_1777(g30672,g16401,g30489);
  nor NOR2_1778(g30673,g16402,g30490);
  nor NOR2_1779(g30674,g16414,g30492);
  nor NOR2_1780(g30675,g16416,g30495);
  nor NOR2_1781(g30676,g16419,g30496);
  nor NOR2_1782(g30677,g16421,g30499);
  nor NOR2_1783(g30678,g16427,g30502);
  nor NOR2_1784(g30679,g16429,g30504);
  nor NOR2_1785(g30680,g16443,g30327);
  nor NOR2_1786(g30681,g16448,g30330);
  nor NOR2_1787(g30682,g16450,g30333);
  nor NOR2_1788(g30683,g16453,g30334);
  nor NOR2_1789(g30684,g16455,g30337);
  nor NOR3_419(g30685,g29992,g30000,g30372);
  nor NOR2_1790(g30686,g16461,g30340);
  nor NOR2_1791(g30687,g13479,g30345);
  nor NOR2_1792(g30688,g13484,g30348);
  nor NOR2_1793(g30689,g13486,g30351);
  nor NOR2_1794(g30690,g13489,g30352);
  nor NOR2_1795(g30691,g13491,g30355);
  nor NOR2_1796(g30692,g13498,g30361);
  nor NOR2_1797(g30693,g13503,g30364);
  nor NOR2_1798(g30694,g13505,g30367);
  nor NOR2_1799(g30695,g13515,g30374);
  nor NOR2_1800(g30699,g13914,g30387);
  nor NOR2_1801(g30700,g13952,g30388);
  nor NOR2_1802(g30701,g13970,g30389);
  nor NOR2_1803(g30702,g14006,g30390);
  nor NOR2_1804(g30703,g14022,g30391);
  nor NOR2_1805(g30704,g14040,g30392);
  nor NOR2_1806(g30705,g14097,g30393);
  nor NOR2_1807(g30706,g14113,g30394);
  nor NOR2_1808(g30707,g14131,g30395);
  nor NOR2_1809(g30708,g14212,g30396);
  nor NOR2_1810(g30709,g14228,g30397);
  nor NOR2_1811(g30780,g30625,g22387);
  nor NOR2_1812(g30783,g30618,g22387);
  nor NOR2_1813(g30785,g30618,g22387);
  nor NOR2_1814(g30786,g30625,g22387);
  nor NOR2_1815(g30787,g30594,g22387);
  nor NOR2_1816(g30788,g30602,g22387);
  nor NOR2_1817(g30789,g30575,g22387);
  nor NOR2_1818(g30790,g30575,g22387);
  nor NOR2_1819(g30796,g16069,g30696);
  nor NOR2_1820(g30798,g16134,g30697);
  nor NOR2_1821(g30801,g16237,g30698);
  nor NOR2_1822(g30929,g30728,g30736);
  nor NOR2_1823(g30930,g30735,g30744);
  nor NOR2_1824(g30931,g30743,g30750);
  nor NOR2_1825(g30932,g30754,g30757);
  nor NOR2_1826(g30933,g30755,g30758);
  nor NOR2_1827(g30934,g30759,g30761);
  nor NOR2_1828(g30935,g30760,g30762);
  nor NOR2_1829(g30936,g30763,g30764);
  nor NOR2_1830(g30954,g30916,g30944);
  nor NOR2_1831(g30955,g30918,g30945);
  nor NOR2_1832(g30956,g30919,g30946);
  nor NOR2_1833(g30957,g30920,g30947);
  nor NOR2_1834(g30958,g30922,g30948);
  nor NOR2_1835(g30959,g30923,g30949);
  nor NOR2_1836(g30960,g30924,g30950);
  nor NOR2_1837(g30961,g30925,g30951);
  nor NOR3_420(g30970,g30917,g30921,g30953);

endmodule
